module load_packet #(
    parameter WIDTH         = 30,
    parameter NUM_PACKET    = 13910,
    parameter NUM_PIC       = 100
)
(
    input                   clk,
    input                   reset_n,
    input                   start,
    input                   ren2in_buf,
    input                   tick,
    input                   packet_out_valid,
    input       [7:0]       packet_out,
    input       [2:0]       grid_state,
    
    output                  input_buffer_empty,
    output                  complete,
    output      [2:0]       state,
    output      [249:0]     spike_out, //dữ liệu ra để ghi vào file txt
    output      [WIDTH-1:0] packet_in, //
    output      [31:0]      num_pack  // 
);
    localparam  [2:0]   IDLE        = 3'b000;
    localparam  [2:0]   LOAD	    = 3'b001;
    localparam  [2:0]   COMPUTE     = 3'b010;
    localparam  [2:0]   WAIT_END    = 3'b100;
    
    reg [WIDTH-1:0]     mem     [0:NUM_PACKET-1];
    reg [9:0]           num_pic [0:NUM_PIC-1];
    reg [31:0]          ptr_packet_reg, ptr_packet_next;
    reg [31:0]          ptr_pic_reg, ptr_pic_next;
    reg [249:0]         compute_out_reg, compute_out_next;
    reg [WIDTH-1:0]     packet_reg, packet_next;
    reg [9:0]           num_line_reg, num_line_next;
    reg [2:0]           state_reg, state_next;
    reg                 complete_reg, complete_next;
    reg [249:0]         spike_reg, spike_next;
    reg                 i_buff_empty_reg, i_buff_empty_next;

    always @(posedge clk or negedge reset_n ) begin
        if (!reset_n) begin
            ptr_packet_reg  <= 0;
            ptr_pic_reg     <= 0;
            state_reg       <= IDLE;
            num_line_reg    <= 0;
            complete_reg    <= 0;
            // mem[0] <= 30'b000000000000000000110010110000
            // ;mem[1] <= 30'b000000000000000000110011000000
            // ;mem[2] <= 30'b000000000000000000110011010000
            // ;mem[3] <= 30'b000000000000000000111001100000
            // ;mem[4] <= 30'b000000000000000000111001110000
            // ;mem[5] <= 30'b000000000000000000111010000000
            // ;mem[6] <= 30'b000000000000000000111010010000
            // ;mem[7] <= 30'b000000000000000000111010100000
            // ;mem[8] <= 30'b000000000000000000111010110000
            // ;mem[9] <= 30'b000000000000000000111011000000
            // ;mem[10] <= 30'b000000000000000000111011010000
            // ;mem[11] <= 30'b000000000000000000111011100000
            // ;mem[12] <= 30'b000000000000000000111011110000
            // ;mem[13] <= 30'b000000000000000000111100000000
            // ;mem[14] <= 30'b000000000000000000111100010000
            // ;mem[15] <= 30'b000000000000000000111100100000
            // ;mem[16] <= 30'b000000000000000000111100110000
            // ;mem[17] <= 30'b000000000000000000111101000000
            // ;mem[18] <= 30'b000000001000000000000110110000
            // ;mem[19] <= 30'b000000001000000000000111000000
            // ;mem[20] <= 30'b000000001000000000000111010000
            // ;mem[21] <= 30'b000000001000000000001101100000
            // ;mem[22] <= 30'b000000001000000000001101110000
            // ;mem[23] <= 30'b000000001000000000001110000000
            // ;mem[24] <= 30'b000000001000000000001110010000
            // ;mem[25] <= 30'b000000001000000000001110100000
            // ;mem[26] <= 30'b000000001000000000001110110000
            // ;mem[27] <= 30'b000000001000000000001111000000
            // ;mem[28] <= 30'b000000001000000000001111010000
            // ;mem[29] <= 30'b000000001000000000001111100000
            // ;mem[30] <= 30'b000000001000000000001111110000
            // ;mem[31] <= 30'b000000001000000000010000000000
            // ;mem[32] <= 30'b000000001000000000010000010000
            // ;mem[33] <= 30'b000000001000000000010000100000
            // ;mem[34] <= 30'b000000001000000000010000110000
            // ;mem[35] <= 30'b000000001000000000010001000000
            // ;mem[36] <= 30'b000000001000000000010101100000
            // ;mem[37] <= 30'b000000001000000000010101110000
            // ;mem[38] <= 30'b000000001000000000010110000000
            // ;mem[39] <= 30'b000000001000000000010110010000
            // ;mem[40] <= 30'b000000001000000000010110100000
            // ;mem[41] <= 30'b000000001000000000010110110000
            // ;mem[42] <= 30'b000000001000000000010111000000
            // ;mem[43] <= 30'b000000001000000000010111010000
            // ;mem[44] <= 30'b000000001000000000010111100000
            // ;mem[45] <= 30'b000000001000000000010111110000
            // ;mem[46] <= 30'b000000001000000000011000000000
            // ;mem[47] <= 30'b000000001000000000011000010000
            // ;mem[48] <= 30'b000000001000000000011110110000
            // ;mem[49] <= 30'b000000001000000000011111000000
            // ;mem[50] <= 30'b000000001000000000100101110000
            // ;mem[51] <= 30'b000000001000000000100110000000
            // ;mem[52] <= 30'b000000001000000000101100100000
            // ;mem[53] <= 30'b000000001000000000101100110000
            // ;mem[54] <= 30'b000000001000000000110011010000
            // ;mem[55] <= 30'b000000001000000000110011100000
            // ;mem[56] <= 30'b000000001000000000110011110000
            // ;mem[57] <= 30'b000000001000000000111010010000
            // ;mem[58] <= 30'b000000001000000000111010100000
            // ;mem[59] <= 30'b000000010000000000000000100000
            // ;mem[60] <= 30'b000000010000000000000000110000
            // ;mem[61] <= 30'b000000010000000000000111010000
            // ;mem[62] <= 30'b000000010000000000000111100000
            // ;mem[63] <= 30'b000000010000000000000111110000
            // ;mem[64] <= 30'b000000010000000000001110010000
            // ;mem[65] <= 30'b000000010000000000001110100000
            // ;mem[66] <= 30'b000000010000000000010101000000
            // ;mem[67] <= 30'b000000010000000000010101010000
            // ;mem[68] <= 30'b000000010000000000010101100000
            // ;mem[69] <= 30'b000000010000000000011100000000
            // ;mem[70] <= 30'b000000010000000000011100010000
            // ;mem[71] <= 30'b000000010000000000100011000000
            // ;mem[72] <= 30'b000000010000000000100011010000
            // ;mem[73] <= 30'b000000010000000000101001110000
            // ;mem[74] <= 30'b000000010000000000101010000000
            // ;mem[75] <= 30'b000000010000000000110000100000
            // ;mem[76] <= 30'b000000010000000000110000110000
            // ;mem[77] <= 30'b000000010000000000110001000000
            // ;mem[78] <= 30'b000000010000000000110111010000
            // ;mem[79] <= 30'b000000010000000000110111100000
            // ;mem[80] <= 30'b000000010000000000110111110000
            // ;mem[81] <= 30'b000000010000000000111110010000
            // ;mem[82] <= 30'b000000010000000000111110100000
            // ;mem[83] <= 30'b000000000000000001000100100000
            // ;mem[84] <= 30'b000000000000000001000100110000
            // ;mem[85] <= 30'b000000000000000001000101000000
            // ;mem[86] <= 30'b000000000000000001001011010000
            // ;mem[87] <= 30'b000000000000000001001011100000
            // ;mem[88] <= 30'b000000000000000001001011110000
            // ;mem[89] <= 30'b000000000000000001010010010000
            // ;mem[90] <= 30'b000000000000000001010010100000
            // ;mem[91] <= 30'b000000000000000001011001000000
            // ;mem[92] <= 30'b000000000000000001011001010000
            // ;mem[93] <= 30'b000000000000000001011111110000
            // ;mem[94] <= 30'b000000000000000001100000000000
            // ;mem[95] <= 30'b000000000000000001100000010000
            // ;mem[96] <= 30'b000000000000000001100110110000
            // ;mem[97] <= 30'b000000000000000001100111000000
            // ;mem[98] <= 30'b000000000000000001100111010000
            // ;mem[99] <= 30'b000000000000000001101101110000
            // ;mem[100] <= 30'b000000000000000001101110000000
            // ;mem[101] <= 30'b000000000000000001101110010000
            // ;mem[102] <= 30'b000000000000000001110100110000
            // ;mem[103] <= 30'b000000000000000001110101000000
            // ;mem[104] <= 30'b000000000000000000011000000000
            // ;mem[105] <= 30'b000000000000000000011000010000
            // ;mem[106] <= 30'b000000000000000000011000100000
            // ;mem[107] <= 30'b000000000000000000011000110000
            // ;mem[108] <= 30'b000000000000000000011110010000
            // ;mem[109] <= 30'b000000000000000000011110100000
            // ;mem[110] <= 30'b000000000000000000011110110000
            // ;mem[111] <= 30'b000000000000000000011111000000
            // ;mem[112] <= 30'b000000000000000000011111010000
            // ;mem[113] <= 30'b000000000000000000011111100000
            // ;mem[114] <= 30'b000000000000000000011111110000
            // ;mem[115] <= 30'b000000000000000000100000000000
            // ;mem[116] <= 30'b000000000000000000100101000000
            // ;mem[117] <= 30'b000000000000000000100101010000
            // ;mem[118] <= 30'b000000000000000000100101100000
            // ;mem[119] <= 30'b000000000000000000100101110000
            // ;mem[120] <= 30'b000000000000000000100110000000
            // ;mem[121] <= 30'b000000000000000000100110010000
            // ;mem[122] <= 30'b000000000000000000100110100000
            // ;mem[123] <= 30'b000000000000000000100110110000
            // ;mem[124] <= 30'b000000000000000000100111000000
            // ;mem[125] <= 30'b000000000000000000101100000000
            // ;mem[126] <= 30'b000000000000000000101100010000
            // ;mem[127] <= 30'b000000000000000000101100100000
            // ;mem[128] <= 30'b000000000000000000101101110000
            // ;mem[129] <= 30'b000000000000000000101110000000
            // ;mem[130] <= 30'b000000000000000000101110010000
            // ;mem[131] <= 30'b000000000000000000110011000000
            // ;mem[132] <= 30'b000000000000000000110011010000
            // ;mem[133] <= 30'b000000000000000000110100110000
            // ;mem[134] <= 30'b000000000000000000110101000000
            // ;mem[135] <= 30'b000000000000000000111011100000
            // ;mem[136] <= 30'b000000000000000000111011110000
            // ;mem[137] <= 30'b000000000000000000111100000000
            // ;mem[138] <= 30'b000000001000000000000000000000
            // ;mem[139] <= 30'b000000001000000000000000010000
            // ;mem[140] <= 30'b000000001000000000000000100000
            // ;mem[141] <= 30'b000000001000000000000001110000
            // ;mem[142] <= 30'b000000001000000000000010000000
            // ;mem[143] <= 30'b000000001000000000000010010000
            // ;mem[144] <= 30'b000000001000000000000111000000
            // ;mem[145] <= 30'b000000001000000000000111010000
            // ;mem[146] <= 30'b000000001000000000001000110000
            // ;mem[147] <= 30'b000000001000000000001001000000
            // ;mem[148] <= 30'b000000001000000000001111100000
            // ;mem[149] <= 30'b000000001000000000001111110000
            // ;mem[150] <= 30'b000000001000000000010000000000
            // ;mem[151] <= 30'b000000001000000000010110100000
            // ;mem[152] <= 30'b000000001000000000010110110000
            // ;mem[153] <= 30'b000000001000000000010111000000
            // ;mem[154] <= 30'b000000001000000000011101010000
            // ;mem[155] <= 30'b000000001000000000011101100000
            // ;mem[156] <= 30'b000000001000000000011101110000
            // ;mem[157] <= 30'b000000001000000000100100000000
            // ;mem[158] <= 30'b000000001000000000100100010000
            // ;mem[159] <= 30'b000000001000000000100100100000
            // ;mem[160] <= 30'b000000001000000000100100110000
            // ;mem[161] <= 30'b000000001000000000101010110000
            // ;mem[162] <= 30'b000000001000000000101011000000
            // ;mem[163] <= 30'b000000001000000000101011010000
            // ;mem[164] <= 30'b000000001000000000101011100000
            // ;mem[165] <= 30'b000000001000000000110001110000
            // ;mem[166] <= 30'b000000001000000000110010000000
            // ;mem[167] <= 30'b000000001000000000110010010000
            // ;mem[168] <= 30'b000000001000000000111000100000
            // ;mem[169] <= 30'b000000001000000000111000110000
            // ;mem[170] <= 30'b000000001000000000111001000000
            // ;mem[171] <= 30'b000000001000000000111001010000
            // ;mem[172] <= 30'b000000001000000000111111100000
            // ;mem[173] <= 30'b000000001000000000111111110000
            // ;mem[174] <= 30'b000000010000000000000101110000
            // ;mem[175] <= 30'b000000010000000000000110000000
            // ;mem[176] <= 30'b000000010000000000000110010000
            // ;mem[177] <= 30'b000000010000000000001100100000
            // ;mem[178] <= 30'b000000010000000000001100110000
            // ;mem[179] <= 30'b000000010000000000001101000000
            // ;mem[180] <= 30'b000000010000000000001101010000
            // ;mem[181] <= 30'b000000010000000000010011100000
            // ;mem[182] <= 30'b000000010000000000010011110000
            // ;mem[183] <= 30'b000000010000000000010100000000
            // ;mem[184] <= 30'b000000010000000000011010010000
            // ;mem[185] <= 30'b000000010000000000011010100000
            // ;mem[186] <= 30'b000000010000000000011010110000
            // ;mem[187] <= 30'b000000010000000000011011000000
            // ;mem[188] <= 30'b000000010000000000100001000000
            // ;mem[189] <= 30'b000000010000000000100001010000
            // ;mem[190] <= 30'b000000010000000000100001100000
            // ;mem[191] <= 30'b000000010000000000100001110000
            // ;mem[192] <= 30'b000000010000000000101000000000
            // ;mem[193] <= 30'b000000010000000000101000010000
            // ;mem[194] <= 30'b000000010000000000101000100000
            // ;mem[195] <= 30'b000000010000000000101111000000
            // ;mem[196] <= 30'b000000010000000000101111010000
            // ;mem[197] <= 30'b000000010000000000101111100000
            // ;mem[198] <= 30'b000000010000000000110010100000
            // ;mem[199] <= 30'b000000010000000000110010110000
            // ;mem[200] <= 30'b000000010000000000110011000000
            // ;mem[201] <= 30'b000000010000000000110011010000
            // ;mem[202] <= 30'b000000010000000000110110000000
            // ;mem[203] <= 30'b000000010000000000110110010000
            // ;mem[204] <= 30'b000000010000000000110110100000
            // ;mem[205] <= 30'b000000010000000000110110110000
            // ;mem[206] <= 30'b000000010000000000110111000000
            // ;mem[207] <= 30'b000000010000000000110111010000
            // ;mem[208] <= 30'b000000010000000000110111100000
            // ;mem[209] <= 30'b000000010000000000110111110000
            // ;mem[210] <= 30'b000000010000000000111000000000
            // ;mem[211] <= 30'b000000010000000000111000010000
            // ;mem[212] <= 30'b000000010000000000111000100000
            // ;mem[213] <= 30'b000000010000000000111000110000
            // ;mem[214] <= 30'b000000010000000000111001000000
            // ;mem[215] <= 30'b000000010000000000111001010000
            // ;mem[216] <= 30'b000000010000000000111001100000
            // ;mem[217] <= 30'b000000010000000000111001110000
            // ;mem[218] <= 30'b000000010000000000111010000000
            // ;mem[219] <= 30'b000000010000000000111010010000
            // ;mem[220] <= 30'b000000010000000000111101000000
            // ;mem[221] <= 30'b000000010000000000111101010000
            // ;mem[222] <= 30'b000000010000000000111101100000
            // ;mem[223] <= 30'b000000010000000000111101110000
            // ;mem[224] <= 30'b000000010000000000111110000000
            // ;mem[225] <= 30'b000000010000000000111110010000
            // ;mem[226] <= 30'b000000010000000000111110100000
            // ;mem[227] <= 30'b000000010000000000111110110000
            // ;mem[228] <= 30'b000000010000000000111111000000
            // ;mem[229] <= 30'b000000010000000000111111010000
            // ;mem[230] <= 30'b000000010000000000111111100000
            // ;mem[231] <= 30'b000000010000000000111111110000
            // ;mem[232] <= 30'b000000000000000001000011000000
            // ;mem[233] <= 30'b000000000000000001000011010000
            // ;mem[234] <= 30'b000000000000000001000011100000
            // ;mem[235] <= 30'b000000000000000001000110100000
            // ;mem[236] <= 30'b000000000000000001000110110000
            // ;mem[237] <= 30'b000000000000000001000111000000
            // ;mem[238] <= 30'b000000000000000001000111010000
            // ;mem[239] <= 30'b000000000000000001001010000000
            // ;mem[240] <= 30'b000000000000000001001010010000
            // ;mem[241] <= 30'b000000000000000001001010100000
            // ;mem[242] <= 30'b000000000000000001001010110000
            // ;mem[243] <= 30'b000000000000000001001011000000
            // ;mem[244] <= 30'b000000000000000001001011010000
            // ;mem[245] <= 30'b000000000000000001001011100000
            // ;mem[246] <= 30'b000000000000000001001011110000
            // ;mem[247] <= 30'b000000000000000001001100000000
            // ;mem[248] <= 30'b000000000000000001001100010000
            // ;mem[249] <= 30'b000000000000000001001100100000
            // ;mem[250] <= 30'b000000000000000001001100110000
            // ;mem[251] <= 30'b000000000000000001001101000000
            // ;mem[252] <= 30'b000000000000000001001101010000
            // ;mem[253] <= 30'b000000000000000001001101100000
            // ;mem[254] <= 30'b000000000000000001001101110000
            // ;mem[255] <= 30'b000000000000000001001110000000
            // ;mem[256] <= 30'b000000000000000001001110010000
            // ;mem[257] <= 30'b000000000000000001010001000000
            // ;mem[258] <= 30'b000000000000000001010001010000
            // ;mem[259] <= 30'b000000000000000001010001100000
            // ;mem[260] <= 30'b000000000000000001010001110000
            // ;mem[261] <= 30'b000000000000000001010010000000
            // ;mem[262] <= 30'b000000000000000001010010010000
            // ;mem[263] <= 30'b000000000000000001010010100000
            // ;mem[264] <= 30'b000000000000000001010010110000
            // ;mem[265] <= 30'b000000000000000001010011000000
            // ;mem[266] <= 30'b000000000000000001010011010000
            // ;mem[267] <= 30'b000000000000000001010011100000
            // ;mem[268] <= 30'b000000000000000001010011110000
            // ;mem[269] <= 30'b000000000000000001010100000000
            // ;mem[270] <= 30'b000000000000000001010100010000
            // ;mem[271] <= 30'b000000000000000001010100100000
            // ;mem[272] <= 30'b000000000000000001010100110000
            // ;mem[273] <= 30'b000000000000000001011001010000
            // ;mem[274] <= 30'b000000000000000001011001100000
            // ;mem[275] <= 30'b000000000000000001011001110000
            // ;mem[276] <= 30'b000000000000000001011010000000
            // ;mem[277] <= 30'b000000000000000001011010010000
            // ;mem[278] <= 30'b000000000000000000100000010000
            // ;mem[279] <= 30'b000000000000000000100111010000
            // ;mem[280] <= 30'b000000000000000000101110000000
            // ;mem[281] <= 30'b000000000000000000101110010000
            // ;mem[282] <= 30'b000000000000000000110101000000
            // ;mem[283] <= 30'b000000000000000000110101010000
            // ;mem[284] <= 30'b000000000000000000111100000000
            // ;mem[285] <= 30'b000000001000000000000010000000
            // ;mem[286] <= 30'b000000001000000000000010010000
            // ;mem[287] <= 30'b000000001000000000001001000000
            // ;mem[288] <= 30'b000000001000000000001001010000
            // ;mem[289] <= 30'b000000001000000000010000000000
            // ;mem[290] <= 30'b000000001000000000010110110000
            // ;mem[291] <= 30'b000000001000000000010111000000
            // ;mem[292] <= 30'b000000001000000000011101110000
            // ;mem[293] <= 30'b000000001000000000011110000000
            // ;mem[294] <= 30'b000000001000000000100100110000
            // ;mem[295] <= 30'b000000001000000000100101000000
            // ;mem[296] <= 30'b000000001000000000101011100000
            // ;mem[297] <= 30'b000000001000000000101011110000
            // ;mem[298] <= 30'b000000001000000000110010100000
            // ;mem[299] <= 30'b000000001000000000110010110000
            // ;mem[300] <= 30'b000000001000000000111001100000
            // ;mem[301] <= 30'b000000001000000000111001110000
            // ;mem[302] <= 30'b000000010000000000000110100000
            // ;mem[303] <= 30'b000000010000000000000110110000
            // ;mem[304] <= 30'b000000010000000000001101100000
            // ;mem[305] <= 30'b000000010000000000001101110000
            // ;mem[306] <= 30'b000000010000000000010100010000
            // ;mem[307] <= 30'b000000010000000000010100100000
            // ;mem[308] <= 30'b000000010000000000011011010000
            // ;mem[309] <= 30'b000000010000000000011011100000
            // ;mem[310] <= 30'b000000010000000000100010010000
            // ;mem[311] <= 30'b000000010000000000100010100000
            // ;mem[312] <= 30'b000000010000000000101001000000
            // ;mem[313] <= 30'b000000010000000000101001010000
            // ;mem[314] <= 30'b000000010000000000101001100000
            // ;mem[315] <= 30'b000000010000000000110000000000
            // ;mem[316] <= 30'b000000010000000000110000010000
            // ;mem[317] <= 30'b000000010000000000110111000000
            // ;mem[318] <= 30'b000000010000000000110111010000
            // ;mem[319] <= 30'b000000010000000000111101110000
            // ;mem[320] <= 30'b000000010000000000111110000000
            // ;mem[321] <= 30'b000000010000000000111110010000
            // ;mem[322] <= 30'b000000000000000001000100000000
            // ;mem[323] <= 30'b000000000000000001000100010000
            // ;mem[324] <= 30'b000000000000000001001011000000
            // ;mem[325] <= 30'b000000000000000001001011010000
            // ;mem[326] <= 30'b000000000000000001010001110000
            // ;mem[327] <= 30'b000000000000000001010010000000
            // ;mem[328] <= 30'b000000000000000001010010010000
            // ;mem[329] <= 30'b000000000000000001011000110000
            // ;mem[330] <= 30'b000000000000000001011001000000
            // ;mem[331] <= 30'b000000000000000001011111110000
            // ;mem[332] <= 30'b000000000000000001100000000000
            // ;mem[333] <= 30'b000000000000000000011111010000
            // ;mem[334] <= 30'b000000000000000000011111100000
            // ;mem[335] <= 30'b000000000000000000011111110000
            // ;mem[336] <= 30'b000000000000000000100110010000
            // ;mem[337] <= 30'b000000000000000000100110100000
            // ;mem[338] <= 30'b000000000000000000100110110000
            // ;mem[339] <= 30'b000000000000000000101101000000
            // ;mem[340] <= 30'b000000000000000000101101010000
            // ;mem[341] <= 30'b000000000000000000101101100000
            // ;mem[342] <= 30'b000000000000000000101101110000
            // ;mem[343] <= 30'b000000000000000000110011110000
            // ;mem[344] <= 30'b000000000000000000110100000000
            // ;mem[345] <= 30'b000000000000000000110100010000
            // ;mem[346] <= 30'b000000000000000000110100100000
            // ;mem[347] <= 30'b000000000000000000110100110000
            // ;mem[348] <= 30'b000000000000000000110101000000
            // ;mem[349] <= 30'b000000000000000000111010100000
            // ;mem[350] <= 30'b000000000000000000111010110000
            // ;mem[351] <= 30'b000000000000000000111011000000
            // ;mem[352] <= 30'b000000000000000000111011010000
            // ;mem[353] <= 30'b000000000000000000111011100000
            // ;mem[354] <= 30'b000000000000000000111011110000
            // ;mem[355] <= 30'b000000000000000000111100000000
            // ;mem[356] <= 30'b000000000000000000111100010000
            // ;mem[357] <= 30'b000000000000000000111100100000
            // ;mem[358] <= 30'b000000001000000000000001000000
            // ;mem[359] <= 30'b000000001000000000000001010000
            // ;mem[360] <= 30'b000000001000000000000001100000
            // ;mem[361] <= 30'b000000001000000000000001110000
            // ;mem[362] <= 30'b000000001000000000000111110000
            // ;mem[363] <= 30'b000000001000000000001000000000
            // ;mem[364] <= 30'b000000001000000000001000010000
            // ;mem[365] <= 30'b000000001000000000001000100000
            // ;mem[366] <= 30'b000000001000000000001000110000
            // ;mem[367] <= 30'b000000001000000000001001000000
            // ;mem[368] <= 30'b000000001000000000001110100000
            // ;mem[369] <= 30'b000000001000000000001110110000
            // ;mem[370] <= 30'b000000001000000000001111000000
            // ;mem[371] <= 30'b000000001000000000001111010000
            // ;mem[372] <= 30'b000000001000000000001111100000
            // ;mem[373] <= 30'b000000001000000000001111110000
            // ;mem[374] <= 30'b000000001000000000010000000000
            // ;mem[375] <= 30'b000000001000000000010000010000
            // ;mem[376] <= 30'b000000001000000000010000100000
            // ;mem[377] <= 30'b000000001000000000010101010000
            // ;mem[378] <= 30'b000000001000000000010101100000
            // ;mem[379] <= 30'b000000001000000000010101110000
            // ;mem[380] <= 30'b000000001000000000010110000000
            // ;mem[381] <= 30'b000000001000000000010110010000
            // ;mem[382] <= 30'b000000001000000000010110100000
            // ;mem[383] <= 30'b000000001000000000010110110000
            // ;mem[384] <= 30'b000000001000000000010111000000
            // ;mem[385] <= 30'b000000001000000000010111010000
            // ;mem[386] <= 30'b000000001000000000010111100000
            // ;mem[387] <= 30'b000000001000000000010111110000
            // ;mem[388] <= 30'b000000001000000000011100010000
            // ;mem[389] <= 30'b000000001000000000011100100000
            // ;mem[390] <= 30'b000000001000000000011100110000
            // ;mem[391] <= 30'b000000001000000000011101000000
            // ;mem[392] <= 30'b000000001000000000011101010000
            // ;mem[393] <= 30'b000000001000000000011101100000
            // ;mem[394] <= 30'b000000001000000000011110010000
            // ;mem[395] <= 30'b000000001000000000011110100000
            // ;mem[396] <= 30'b000000001000000000011110110000
            // ;mem[397] <= 30'b000000001000000000100011000000
            // ;mem[398] <= 30'b000000001000000000100011010000
            // ;mem[399] <= 30'b000000001000000000100011100000
            // ;mem[400] <= 30'b000000001000000000100011110000
            // ;mem[401] <= 30'b000000001000000000100100000000
            // ;mem[402] <= 30'b000000001000000000100100010000
            // ;mem[403] <= 30'b000000001000000000100101100000
            // ;mem[404] <= 30'b000000001000000000100101110000
            // ;mem[405] <= 30'b000000001000000000100110000000
            // ;mem[406] <= 30'b000000001000000000101010000000
            // ;mem[407] <= 30'b000000001000000000101010010000
            // ;mem[408] <= 30'b000000001000000000101010100000
            // ;mem[409] <= 30'b000000001000000000101010110000
            // ;mem[410] <= 30'b000000001000000000101100110000
            // ;mem[411] <= 30'b000000001000000000101101000000
            // ;mem[412] <= 30'b000000001000000000101101010000
            // ;mem[413] <= 30'b000000001000000000110001000000
            // ;mem[414] <= 30'b000000001000000000110001010000
            // ;mem[415] <= 30'b000000001000000000110001100000
            // ;mem[416] <= 30'b000000001000000000110011110000
            // ;mem[417] <= 30'b000000001000000000110100000000
            // ;mem[418] <= 30'b000000001000000000110100010000
            // ;mem[419] <= 30'b000000001000000000111000000000
            // ;mem[420] <= 30'b000000001000000000111000010000
            // ;mem[421] <= 30'b000000001000000000111010110000
            // ;mem[422] <= 30'b000000001000000000111011000000
            // ;mem[423] <= 30'b000000001000000000111011010000
            // ;mem[424] <= 30'b000000001000000000111011100000
            // ;mem[425] <= 30'b000000001000000000111110110000
            // ;mem[426] <= 30'b000000001000000000111111000000
            // ;mem[427] <= 30'b000000001000000000111111010000
            // ;mem[428] <= 30'b000000010000000000000000110000
            // ;mem[429] <= 30'b000000010000000000000001000000
            // ;mem[430] <= 30'b000000010000000000000001010000
            // ;mem[431] <= 30'b000000010000000000000101000000
            // ;mem[432] <= 30'b000000010000000000000101010000
            // ;mem[433] <= 30'b000000010000000000000101100000
            // ;mem[434] <= 30'b000000010000000000000111110000
            // ;mem[435] <= 30'b000000010000000000001000000000
            // ;mem[436] <= 30'b000000010000000000001000010000
            // ;mem[437] <= 30'b000000010000000000001100000000
            // ;mem[438] <= 30'b000000010000000000001100010000
            // ;mem[439] <= 30'b000000010000000000001110110000
            // ;mem[440] <= 30'b000000010000000000001111000000
            // ;mem[441] <= 30'b000000010000000000001111010000
            // ;mem[442] <= 30'b000000010000000000001111100000
            // ;mem[443] <= 30'b000000010000000000010010110000
            // ;mem[444] <= 30'b000000010000000000010011000000
            // ;mem[445] <= 30'b000000010000000000010011010000
            // ;mem[446] <= 30'b000000010000000000010101110000
            // ;mem[447] <= 30'b000000010000000000010110000000
            // ;mem[448] <= 30'b000000010000000000010110010000
            // ;mem[449] <= 30'b000000010000000000011001110000
            // ;mem[450] <= 30'b000000010000000000011010000000
            // ;mem[451] <= 30'b000000010000000000011010010000
            // ;mem[452] <= 30'b000000010000000000011100100000
            // ;mem[453] <= 30'b000000010000000000011100110000
            // ;mem[454] <= 30'b000000010000000000011101000000
            // ;mem[455] <= 30'b000000010000000000011101010000
            // ;mem[456] <= 30'b000000010000000000100000110000
            // ;mem[457] <= 30'b000000010000000000100001000000
            // ;mem[458] <= 30'b000000010000000000100001010000
            // ;mem[459] <= 30'b000000010000000000100011000000
            // ;mem[460] <= 30'b000000010000000000100011010000
            // ;mem[461] <= 30'b000000010000000000100011100000
            // ;mem[462] <= 30'b000000010000000000100011110000
            // ;mem[463] <= 30'b000000010000000000100100000000
            // ;mem[464] <= 30'b000000010000000000100111110000
            // ;mem[465] <= 30'b000000010000000000101000000000
            // ;mem[466] <= 30'b000000010000000000101000010000
            // ;mem[467] <= 30'b000000010000000000101001110000
            // ;mem[468] <= 30'b000000010000000000101010000000
            // ;mem[469] <= 30'b000000010000000000101010010000
            // ;mem[470] <= 30'b000000010000000000101010100000
            // ;mem[471] <= 30'b000000010000000000101010110000
            // ;mem[472] <= 30'b000000010000000000101011000000
            // ;mem[473] <= 30'b000000010000000000101110110000
            // ;mem[474] <= 30'b000000010000000000101111000000
            // ;mem[475] <= 30'b000000010000000000101111010000
            // ;mem[476] <= 30'b000000010000000000110000000000
            // ;mem[477] <= 30'b000000010000000000110000010000
            // ;mem[478] <= 30'b000000010000000000110000100000
            // ;mem[479] <= 30'b000000010000000000110000110000
            // ;mem[480] <= 30'b000000010000000000110001000000
            // ;mem[481] <= 30'b000000010000000000110001010000
            // ;mem[482] <= 30'b000000010000000000110001100000
            // ;mem[483] <= 30'b000000010000000000110001110000
            // ;mem[484] <= 30'b000000010000000000110110000000
            // ;mem[485] <= 30'b000000010000000000110110010000
            // ;mem[486] <= 30'b000000010000000000110110100000
            // ;mem[487] <= 30'b000000010000000000110110110000
            // ;mem[488] <= 30'b000000010000000000110111000000
            // ;mem[489] <= 30'b000000010000000000110111010000
            // ;mem[490] <= 30'b000000010000000000110111100000
            // ;mem[491] <= 30'b000000010000000000110111110000
            // ;mem[492] <= 30'b000000010000000000111000000000
            // ;mem[493] <= 30'b000000010000000000111000010000
            // ;mem[494] <= 30'b000000010000000000111000100000
            // ;mem[495] <= 30'b000000010000000000111000110000
            // ;mem[496] <= 30'b000000010000000000111101000000
            // ;mem[497] <= 30'b000000010000000000111101010000
            // ;mem[498] <= 30'b000000010000000000111101100000
            // ;mem[499] <= 30'b000000010000000000111101110000
            // ;mem[500] <= 30'b000000010000000000111110000000
            // ;mem[501] <= 30'b000000010000000000111110010000
            // ;mem[502] <= 30'b000000010000000000111110100000
            // ;mem[503] <= 30'b000000010000000000111110110000
            // ;mem[504] <= 30'b000000010000000000111111000000
            // ;mem[505] <= 30'b000000010000000000111111010000
            // ;mem[506] <= 30'b000000000000000001000010110000
            // ;mem[507] <= 30'b000000000000000001000011000000
            // ;mem[508] <= 30'b000000000000000001000011010000
            // ;mem[509] <= 30'b000000000000000001000100000000
            // ;mem[510] <= 30'b000000000000000001000100010000
            // ;mem[511] <= 30'b000000000000000001000100100000
            // ;mem[512] <= 30'b000000000000000001000100110000
            // ;mem[513] <= 30'b000000000000000001000101000000
            // ;mem[514] <= 30'b000000000000000001000101010000
            // ;mem[515] <= 30'b000000000000000001000101100000
            // ;mem[516] <= 30'b000000000000000001000101110000
            // ;mem[517] <= 30'b000000000000000001001010000000
            // ;mem[518] <= 30'b000000000000000001001010010000
            // ;mem[519] <= 30'b000000000000000001001010100000
            // ;mem[520] <= 30'b000000000000000001001010110000
            // ;mem[521] <= 30'b000000000000000001001011000000
            // ;mem[522] <= 30'b000000000000000001001011010000
            // ;mem[523] <= 30'b000000000000000001001011100000
            // ;mem[524] <= 30'b000000000000000001001011110000
            // ;mem[525] <= 30'b000000000000000001001100000000
            // ;mem[526] <= 30'b000000000000000001001100010000
            // ;mem[527] <= 30'b000000000000000001001100100000
            // ;mem[528] <= 30'b000000000000000001001100110000
            // ;mem[529] <= 30'b000000000000000001010001000000
            // ;mem[530] <= 30'b000000000000000001010001010000
            // ;mem[531] <= 30'b000000000000000001010001100000
            // ;mem[532] <= 30'b000000000000000001010001110000
            // ;mem[533] <= 30'b000000000000000001010010000000
            // ;mem[534] <= 30'b000000000000000001010010010000
            // ;mem[535] <= 30'b000000000000000001010010100000
            // ;mem[536] <= 30'b000000000000000001010010110000
            // ;mem[537] <= 30'b000000000000000001010011000000
            // ;mem[538] <= 30'b000000000000000001010011010000
            // ;mem[539] <= 30'b000000000000000001011000010000
            // ;mem[540] <= 30'b000000000000000001011000100000
            // ;mem[541] <= 30'b000000000000000001011000110000
            // ;mem[542] <= 30'b000000000000000001011001000000
            // ;mem[543] <= 30'b000000000000000001011001010000
            // ;mem[544] <= 30'b000000000000000001011001100000
            // ;mem[545] <= 30'b000000000000000001011001110000
            // ;mem[546] <= 30'b000000000000000001011111110000
            // ;mem[547] <= 30'b000000000000000001100000000000
            // ;mem[548] <= 30'b000000000000000001100000010000;
            // num_pic[0] <= 10'h68;
            // num_pic[1] <= 10'hae;
            // num_pic[2] <= 10'h37;
            // num_pic[3] <= 10'hd8;
            //All packet
                num_pic[0] <= 10'h68
                ;num_pic[1] <= 10'hae
                ;num_pic[2] <= 10'h37
                ;num_pic[3] <= 10'hd8
                ;num_pic[4] <= 10'h6a
                ;num_pic[5] <= 10'h50
                ;num_pic[6] <= 10'h88
                ;num_pic[7] <= 10'h77
                ;num_pic[8] <= 10'hbb
                ;num_pic[9] <= 10'hbe
                ;num_pic[10] <= 10'hb4
                ;num_pic[11] <= 10'ha5
                ;num_pic[12] <= 10'h83
                ;num_pic[13] <= 10'ha9
                ;num_pic[14] <= 10'h65
                ;num_pic[15] <= 10'h71
                ;num_pic[16] <= 10'h80
                ;num_pic[17] <= 10'h7b
                ;num_pic[18] <= 10'hcd
                ;num_pic[19] <= 10'h52
                ;num_pic[20] <= 10'h9b
                ;num_pic[21] <= 10'h8a
                ;num_pic[22] <= 10'h82
                ;num_pic[23] <= 10'h78
                ;num_pic[24] <= 10'h4b
                ;num_pic[25] <= 10'h134
                ;num_pic[26] <= 10'h51
                ;num_pic[27] <= 10'h81
                ;num_pic[28] <= 10'hc9
                ;num_pic[29] <= 10'h44
                ;num_pic[30] <= 10'h98
                ;num_pic[31] <= 10'h3c
                ;num_pic[32] <= 10'h93
                ;num_pic[33] <= 10'h8b
                ;num_pic[34] <= 10'h99
                ;num_pic[35] <= 10'hae
                ;num_pic[36] <= 10'h87
                ;num_pic[37] <= 10'h50
                ;num_pic[38] <= 10'h72
                ;num_pic[39] <= 10'h6b
                ;num_pic[40] <= 10'h25
                ;num_pic[41] <= 10'h5b
                ;num_pic[42] <= 10'h8c
                ;num_pic[43] <= 10'h50
                ;num_pic[44] <= 10'h74
                ;num_pic[45] <= 10'h72
                ;num_pic[46] <= 10'h6c
                ;num_pic[47] <= 10'h57
                ;num_pic[48] <= 10'hdb
                ;num_pic[49] <= 10'h80
                ;num_pic[50] <= 10'h7b
                ;num_pic[51] <= 10'hf7
                ;num_pic[52] <= 10'h82
                ;num_pic[53] <= 10'h5e
                ;num_pic[54] <= 10'hd0
                ;num_pic[55] <= 10'ha1
                ;num_pic[56] <= 10'ha3
                ;num_pic[57] <= 10'h39
                ;num_pic[58] <= 10'h94
                ;num_pic[59] <= 10'h3c
                ;num_pic[60] <= 10'h9c
                ;num_pic[61] <= 10'hce
                ;num_pic[62] <= 10'h53
                ;num_pic[63] <= 10'h8c
                ;num_pic[64] <= 10'hb3
                ;num_pic[65] <= 10'h57
                ;num_pic[66] <= 10'h90
                ;num_pic[67] <= 10'h79
                ;num_pic[68] <= 10'he6
                ;num_pic[69] <= 10'hbe
                ;num_pic[70] <= 10'h7e
                ;num_pic[71] <= 10'hfe
                ;num_pic[72] <= 10'h9e
                ;num_pic[73] <= 10'hac
                ;num_pic[74] <= 10'h58
                ;num_pic[75] <= 10'h69
                ;num_pic[76] <= 10'h69
                ;num_pic[77] <= 10'h70
                ;num_pic[78] <= 10'h75
                ;num_pic[79] <= 10'hce
                ;num_pic[80] <= 10'h76
                ;num_pic[81] <= 10'h9f
                ;num_pic[82] <= 10'hbf
                ;num_pic[83] <= 10'h64
                ;num_pic[84] <= 10'h9a
                ;num_pic[85] <= 10'hdb
                ;num_pic[86] <= 10'h8f
                ;num_pic[87] <= 10'h98
                ;num_pic[88] <= 10'ha6
                ;num_pic[89] <= 10'h62
                ;num_pic[90] <= 10'h94
                ;num_pic[91] <= 10'h84
                ;num_pic[92] <= 10'h54
                ;num_pic[93] <= 10'hd6
                ;num_pic[94] <= 10'h82
                ;num_pic[95] <= 10'hea
                ;num_pic[96] <= 10'h44
                ;num_pic[97] <= 10'had
                ;num_pic[98] <= 10'h86
                ;num_pic[99] <= 10'had;
                mem[0] <= 30'b000000000000000000110010110000
                ;mem[1] <= 30'b000000000000000000110011000000
                ;mem[2] <= 30'b000000000000000000110011010000
                ;mem[3] <= 30'b000000000000000000111001100000
                ;mem[4] <= 30'b000000000000000000111001110000
                ;mem[5] <= 30'b000000000000000000111010000000
                ;mem[6] <= 30'b000000000000000000111010010000
                ;mem[7] <= 30'b000000000000000000111010100000
                ;mem[8] <= 30'b000000000000000000111010110000
                ;mem[9] <= 30'b000000000000000000111011000000
                ;mem[10] <= 30'b000000000000000000111011010000
                ;mem[11] <= 30'b000000000000000000111011100000
                ;mem[12] <= 30'b000000000000000000111011110000
                ;mem[13] <= 30'b000000000000000000111100000000
                ;mem[14] <= 30'b000000000000000000111100010000
                ;mem[15] <= 30'b000000000000000000111100100000
                ;mem[16] <= 30'b000000000000000000111100110000
                ;mem[17] <= 30'b000000000000000000111101000000
                ;mem[18] <= 30'b000000001000000000000110110000
                ;mem[19] <= 30'b000000001000000000000111000000
                ;mem[20] <= 30'b000000001000000000000111010000
                ;mem[21] <= 30'b000000001000000000001101100000
                ;mem[22] <= 30'b000000001000000000001101110000
                ;mem[23] <= 30'b000000001000000000001110000000
                ;mem[24] <= 30'b000000001000000000001110010000
                ;mem[25] <= 30'b000000001000000000001110100000
                ;mem[26] <= 30'b000000001000000000001110110000
                ;mem[27] <= 30'b000000001000000000001111000000
                ;mem[28] <= 30'b000000001000000000001111010000
                ;mem[29] <= 30'b000000001000000000001111100000
                ;mem[30] <= 30'b000000001000000000001111110000
                ;mem[31] <= 30'b000000001000000000010000000000
                ;mem[32] <= 30'b000000001000000000010000010000
                ;mem[33] <= 30'b000000001000000000010000100000
                ;mem[34] <= 30'b000000001000000000010000110000
                ;mem[35] <= 30'b000000001000000000010001000000
                ;mem[36] <= 30'b000000001000000000010101100000
                ;mem[37] <= 30'b000000001000000000010101110000
                ;mem[38] <= 30'b000000001000000000010110000000
                ;mem[39] <= 30'b000000001000000000010110010000
                ;mem[40] <= 30'b000000001000000000010110100000
                ;mem[41] <= 30'b000000001000000000010110110000
                ;mem[42] <= 30'b000000001000000000010111000000
                ;mem[43] <= 30'b000000001000000000010111010000
                ;mem[44] <= 30'b000000001000000000010111100000
                ;mem[45] <= 30'b000000001000000000010111110000
                ;mem[46] <= 30'b000000001000000000011000000000
                ;mem[47] <= 30'b000000001000000000011000010000
                ;mem[48] <= 30'b000000001000000000011110110000
                ;mem[49] <= 30'b000000001000000000011111000000
                ;mem[50] <= 30'b000000001000000000100101110000
                ;mem[51] <= 30'b000000001000000000100110000000
                ;mem[52] <= 30'b000000001000000000101100100000
                ;mem[53] <= 30'b000000001000000000101100110000
                ;mem[54] <= 30'b000000001000000000110011010000
                ;mem[55] <= 30'b000000001000000000110011100000
                ;mem[56] <= 30'b000000001000000000110011110000
                ;mem[57] <= 30'b000000001000000000111010010000
                ;mem[58] <= 30'b000000001000000000111010100000
                ;mem[59] <= 30'b000000010000000000000000100000
                ;mem[60] <= 30'b000000010000000000000000110000
                ;mem[61] <= 30'b000000010000000000000111010000
                ;mem[62] <= 30'b000000010000000000000111100000
                ;mem[63] <= 30'b000000010000000000000111110000
                ;mem[64] <= 30'b000000010000000000001110010000
                ;mem[65] <= 30'b000000010000000000001110100000
                ;mem[66] <= 30'b000000010000000000010101000000
                ;mem[67] <= 30'b000000010000000000010101010000
                ;mem[68] <= 30'b000000010000000000010101100000
                ;mem[69] <= 30'b000000010000000000011100000000
                ;mem[70] <= 30'b000000010000000000011100010000
                ;mem[71] <= 30'b000000010000000000100011000000
                ;mem[72] <= 30'b000000010000000000100011010000
                ;mem[73] <= 30'b000000010000000000101001110000
                ;mem[74] <= 30'b000000010000000000101010000000
                ;mem[75] <= 30'b000000010000000000110000100000
                ;mem[76] <= 30'b000000010000000000110000110000
                ;mem[77] <= 30'b000000010000000000110001000000
                ;mem[78] <= 30'b000000010000000000110111010000
                ;mem[79] <= 30'b000000010000000000110111100000
                ;mem[80] <= 30'b000000010000000000110111110000
                ;mem[81] <= 30'b000000010000000000111110010000
                ;mem[82] <= 30'b000000010000000000111110100000
                ;mem[83] <= 30'b000000000000000001000100100000
                ;mem[84] <= 30'b000000000000000001000100110000
                ;mem[85] <= 30'b000000000000000001000101000000
                ;mem[86] <= 30'b000000000000000001001011010000
                ;mem[87] <= 30'b000000000000000001001011100000
                ;mem[88] <= 30'b000000000000000001001011110000
                ;mem[89] <= 30'b000000000000000001010010010000
                ;mem[90] <= 30'b000000000000000001010010100000
                ;mem[91] <= 30'b000000000000000001011001000000
                ;mem[92] <= 30'b000000000000000001011001010000
                ;mem[93] <= 30'b000000000000000001011111110000
                ;mem[94] <= 30'b000000000000000001100000000000
                ;mem[95] <= 30'b000000000000000001100000010000
                ;mem[96] <= 30'b000000000000000001100110110000
                ;mem[97] <= 30'b000000000000000001100111000000
                ;mem[98] <= 30'b000000000000000001100111010000
                ;mem[99] <= 30'b000000000000000001101101110000
                ;mem[100] <= 30'b000000000000000001101110000000
                ;mem[101] <= 30'b000000000000000001101110010000
                ;mem[102] <= 30'b000000000000000001110100110000
                ;mem[103] <= 30'b000000000000000001110101000000
                ;mem[104] <= 30'b000000000000000000011000000000
                ;mem[105] <= 30'b000000000000000000011000010000
                ;mem[106] <= 30'b000000000000000000011000100000
                ;mem[107] <= 30'b000000000000000000011000110000
                ;mem[108] <= 30'b000000000000000000011110010000
                ;mem[109] <= 30'b000000000000000000011110100000
                ;mem[110] <= 30'b000000000000000000011110110000
                ;mem[111] <= 30'b000000000000000000011111000000
                ;mem[112] <= 30'b000000000000000000011111010000
                ;mem[113] <= 30'b000000000000000000011111100000
                ;mem[114] <= 30'b000000000000000000011111110000
                ;mem[115] <= 30'b000000000000000000100000000000
                ;mem[116] <= 30'b000000000000000000100101000000
                ;mem[117] <= 30'b000000000000000000100101010000
                ;mem[118] <= 30'b000000000000000000100101100000
                ;mem[119] <= 30'b000000000000000000100101110000
                ;mem[120] <= 30'b000000000000000000100110000000
                ;mem[121] <= 30'b000000000000000000100110010000
                ;mem[122] <= 30'b000000000000000000100110100000
                ;mem[123] <= 30'b000000000000000000100110110000
                ;mem[124] <= 30'b000000000000000000100111000000
                ;mem[125] <= 30'b000000000000000000101100000000
                ;mem[126] <= 30'b000000000000000000101100010000
                ;mem[127] <= 30'b000000000000000000101100100000
                ;mem[128] <= 30'b000000000000000000101101110000
                ;mem[129] <= 30'b000000000000000000101110000000
                ;mem[130] <= 30'b000000000000000000101110010000
                ;mem[131] <= 30'b000000000000000000110011000000
                ;mem[132] <= 30'b000000000000000000110011010000
                ;mem[133] <= 30'b000000000000000000110100110000
                ;mem[134] <= 30'b000000000000000000110101000000
                ;mem[135] <= 30'b000000000000000000111011100000
                ;mem[136] <= 30'b000000000000000000111011110000
                ;mem[137] <= 30'b000000000000000000111100000000
                ;mem[138] <= 30'b000000001000000000000000000000
                ;mem[139] <= 30'b000000001000000000000000010000
                ;mem[140] <= 30'b000000001000000000000000100000
                ;mem[141] <= 30'b000000001000000000000001110000
                ;mem[142] <= 30'b000000001000000000000010000000
                ;mem[143] <= 30'b000000001000000000000010010000
                ;mem[144] <= 30'b000000001000000000000111000000
                ;mem[145] <= 30'b000000001000000000000111010000
                ;mem[146] <= 30'b000000001000000000001000110000
                ;mem[147] <= 30'b000000001000000000001001000000
                ;mem[148] <= 30'b000000001000000000001111100000
                ;mem[149] <= 30'b000000001000000000001111110000
                ;mem[150] <= 30'b000000001000000000010000000000
                ;mem[151] <= 30'b000000001000000000010110100000
                ;mem[152] <= 30'b000000001000000000010110110000
                ;mem[153] <= 30'b000000001000000000010111000000
                ;mem[154] <= 30'b000000001000000000011101010000
                ;mem[155] <= 30'b000000001000000000011101100000
                ;mem[156] <= 30'b000000001000000000011101110000
                ;mem[157] <= 30'b000000001000000000100100000000
                ;mem[158] <= 30'b000000001000000000100100010000
                ;mem[159] <= 30'b000000001000000000100100100000
                ;mem[160] <= 30'b000000001000000000100100110000
                ;mem[161] <= 30'b000000001000000000101010110000
                ;mem[162] <= 30'b000000001000000000101011000000
                ;mem[163] <= 30'b000000001000000000101011010000
                ;mem[164] <= 30'b000000001000000000101011100000
                ;mem[165] <= 30'b000000001000000000110001110000
                ;mem[166] <= 30'b000000001000000000110010000000
                ;mem[167] <= 30'b000000001000000000110010010000
                ;mem[168] <= 30'b000000001000000000111000100000
                ;mem[169] <= 30'b000000001000000000111000110000
                ;mem[170] <= 30'b000000001000000000111001000000
                ;mem[171] <= 30'b000000001000000000111001010000
                ;mem[172] <= 30'b000000001000000000111111100000
                ;mem[173] <= 30'b000000001000000000111111110000
                ;mem[174] <= 30'b000000010000000000000101110000
                ;mem[175] <= 30'b000000010000000000000110000000
                ;mem[176] <= 30'b000000010000000000000110010000
                ;mem[177] <= 30'b000000010000000000001100100000
                ;mem[178] <= 30'b000000010000000000001100110000
                ;mem[179] <= 30'b000000010000000000001101000000
                ;mem[180] <= 30'b000000010000000000001101010000
                ;mem[181] <= 30'b000000010000000000010011100000
                ;mem[182] <= 30'b000000010000000000010011110000
                ;mem[183] <= 30'b000000010000000000010100000000
                ;mem[184] <= 30'b000000010000000000011010010000
                ;mem[185] <= 30'b000000010000000000011010100000
                ;mem[186] <= 30'b000000010000000000011010110000
                ;mem[187] <= 30'b000000010000000000011011000000
                ;mem[188] <= 30'b000000010000000000100001000000
                ;mem[189] <= 30'b000000010000000000100001010000
                ;mem[190] <= 30'b000000010000000000100001100000
                ;mem[191] <= 30'b000000010000000000100001110000
                ;mem[192] <= 30'b000000010000000000101000000000
                ;mem[193] <= 30'b000000010000000000101000010000
                ;mem[194] <= 30'b000000010000000000101000100000
                ;mem[195] <= 30'b000000010000000000101111000000
                ;mem[196] <= 30'b000000010000000000101111010000
                ;mem[197] <= 30'b000000010000000000101111100000
                ;mem[198] <= 30'b000000010000000000110010100000
                ;mem[199] <= 30'b000000010000000000110010110000
                ;mem[200] <= 30'b000000010000000000110011000000
                ;mem[201] <= 30'b000000010000000000110011010000
                ;mem[202] <= 30'b000000010000000000110110000000
                ;mem[203] <= 30'b000000010000000000110110010000
                ;mem[204] <= 30'b000000010000000000110110100000
                ;mem[205] <= 30'b000000010000000000110110110000
                ;mem[206] <= 30'b000000010000000000110111000000
                ;mem[207] <= 30'b000000010000000000110111010000
                ;mem[208] <= 30'b000000010000000000110111100000
                ;mem[209] <= 30'b000000010000000000110111110000
                ;mem[210] <= 30'b000000010000000000111000000000
                ;mem[211] <= 30'b000000010000000000111000010000
                ;mem[212] <= 30'b000000010000000000111000100000
                ;mem[213] <= 30'b000000010000000000111000110000
                ;mem[214] <= 30'b000000010000000000111001000000
                ;mem[215] <= 30'b000000010000000000111001010000
                ;mem[216] <= 30'b000000010000000000111001100000
                ;mem[217] <= 30'b000000010000000000111001110000
                ;mem[218] <= 30'b000000010000000000111010000000
                ;mem[219] <= 30'b000000010000000000111010010000
                ;mem[220] <= 30'b000000010000000000111101000000
                ;mem[221] <= 30'b000000010000000000111101010000
                ;mem[222] <= 30'b000000010000000000111101100000
                ;mem[223] <= 30'b000000010000000000111101110000
                ;mem[224] <= 30'b000000010000000000111110000000
                ;mem[225] <= 30'b000000010000000000111110010000
                ;mem[226] <= 30'b000000010000000000111110100000
                ;mem[227] <= 30'b000000010000000000111110110000
                ;mem[228] <= 30'b000000010000000000111111000000
                ;mem[229] <= 30'b000000010000000000111111010000
                ;mem[230] <= 30'b000000010000000000111111100000
                ;mem[231] <= 30'b000000010000000000111111110000
                ;mem[232] <= 30'b000000000000000001000011000000
                ;mem[233] <= 30'b000000000000000001000011010000
                ;mem[234] <= 30'b000000000000000001000011100000
                ;mem[235] <= 30'b000000000000000001000110100000
                ;mem[236] <= 30'b000000000000000001000110110000
                ;mem[237] <= 30'b000000000000000001000111000000
                ;mem[238] <= 30'b000000000000000001000111010000
                ;mem[239] <= 30'b000000000000000001001010000000
                ;mem[240] <= 30'b000000000000000001001010010000
                ;mem[241] <= 30'b000000000000000001001010100000
                ;mem[242] <= 30'b000000000000000001001010110000
                ;mem[243] <= 30'b000000000000000001001011000000
                ;mem[244] <= 30'b000000000000000001001011010000
                ;mem[245] <= 30'b000000000000000001001011100000
                ;mem[246] <= 30'b000000000000000001001011110000
                ;mem[247] <= 30'b000000000000000001001100000000
                ;mem[248] <= 30'b000000000000000001001100010000
                ;mem[249] <= 30'b000000000000000001001100100000
                ;mem[250] <= 30'b000000000000000001001100110000
                ;mem[251] <= 30'b000000000000000001001101000000
                ;mem[252] <= 30'b000000000000000001001101010000
                ;mem[253] <= 30'b000000000000000001001101100000
                ;mem[254] <= 30'b000000000000000001001101110000
                ;mem[255] <= 30'b000000000000000001001110000000
                ;mem[256] <= 30'b000000000000000001001110010000
                ;mem[257] <= 30'b000000000000000001010001000000
                ;mem[258] <= 30'b000000000000000001010001010000
                ;mem[259] <= 30'b000000000000000001010001100000
                ;mem[260] <= 30'b000000000000000001010001110000
                ;mem[261] <= 30'b000000000000000001010010000000
                ;mem[262] <= 30'b000000000000000001010010010000
                ;mem[263] <= 30'b000000000000000001010010100000
                ;mem[264] <= 30'b000000000000000001010010110000
                ;mem[265] <= 30'b000000000000000001010011000000
                ;mem[266] <= 30'b000000000000000001010011010000
                ;mem[267] <= 30'b000000000000000001010011100000
                ;mem[268] <= 30'b000000000000000001010011110000
                ;mem[269] <= 30'b000000000000000001010100000000
                ;mem[270] <= 30'b000000000000000001010100010000
                ;mem[271] <= 30'b000000000000000001010100100000
                ;mem[272] <= 30'b000000000000000001010100110000
                ;mem[273] <= 30'b000000000000000001011001010000
                ;mem[274] <= 30'b000000000000000001011001100000
                ;mem[275] <= 30'b000000000000000001011001110000
                ;mem[276] <= 30'b000000000000000001011010000000
                ;mem[277] <= 30'b000000000000000001011010010000
                ;mem[278] <= 30'b000000000000000000100000010000
                ;mem[279] <= 30'b000000000000000000100111010000
                ;mem[280] <= 30'b000000000000000000101110000000
                ;mem[281] <= 30'b000000000000000000101110010000
                ;mem[282] <= 30'b000000000000000000110101000000
                ;mem[283] <= 30'b000000000000000000110101010000
                ;mem[284] <= 30'b000000000000000000111100000000
                ;mem[285] <= 30'b000000001000000000000010000000
                ;mem[286] <= 30'b000000001000000000000010010000
                ;mem[287] <= 30'b000000001000000000001001000000
                ;mem[288] <= 30'b000000001000000000001001010000
                ;mem[289] <= 30'b000000001000000000010000000000
                ;mem[290] <= 30'b000000001000000000010110110000
                ;mem[291] <= 30'b000000001000000000010111000000
                ;mem[292] <= 30'b000000001000000000011101110000
                ;mem[293] <= 30'b000000001000000000011110000000
                ;mem[294] <= 30'b000000001000000000100100110000
                ;mem[295] <= 30'b000000001000000000100101000000
                ;mem[296] <= 30'b000000001000000000101011100000
                ;mem[297] <= 30'b000000001000000000101011110000
                ;mem[298] <= 30'b000000001000000000110010100000
                ;mem[299] <= 30'b000000001000000000110010110000
                ;mem[300] <= 30'b000000001000000000111001100000
                ;mem[301] <= 30'b000000001000000000111001110000
                ;mem[302] <= 30'b000000010000000000000110100000
                ;mem[303] <= 30'b000000010000000000000110110000
                ;mem[304] <= 30'b000000010000000000001101100000
                ;mem[305] <= 30'b000000010000000000001101110000
                ;mem[306] <= 30'b000000010000000000010100010000
                ;mem[307] <= 30'b000000010000000000010100100000
                ;mem[308] <= 30'b000000010000000000011011010000
                ;mem[309] <= 30'b000000010000000000011011100000
                ;mem[310] <= 30'b000000010000000000100010010000
                ;mem[311] <= 30'b000000010000000000100010100000
                ;mem[312] <= 30'b000000010000000000101001000000
                ;mem[313] <= 30'b000000010000000000101001010000
                ;mem[314] <= 30'b000000010000000000101001100000
                ;mem[315] <= 30'b000000010000000000110000000000
                ;mem[316] <= 30'b000000010000000000110000010000
                ;mem[317] <= 30'b000000010000000000110111000000
                ;mem[318] <= 30'b000000010000000000110111010000
                ;mem[319] <= 30'b000000010000000000111101110000
                ;mem[320] <= 30'b000000010000000000111110000000
                ;mem[321] <= 30'b000000010000000000111110010000
                ;mem[322] <= 30'b000000000000000001000100000000
                ;mem[323] <= 30'b000000000000000001000100010000
                ;mem[324] <= 30'b000000000000000001001011000000
                ;mem[325] <= 30'b000000000000000001001011010000
                ;mem[326] <= 30'b000000000000000001010001110000
                ;mem[327] <= 30'b000000000000000001010010000000
                ;mem[328] <= 30'b000000000000000001010010010000
                ;mem[329] <= 30'b000000000000000001011000110000
                ;mem[330] <= 30'b000000000000000001011001000000
                ;mem[331] <= 30'b000000000000000001011111110000
                ;mem[332] <= 30'b000000000000000001100000000000
                ;mem[333] <= 30'b000000000000000000011111010000
                ;mem[334] <= 30'b000000000000000000011111100000
                ;mem[335] <= 30'b000000000000000000011111110000
                ;mem[336] <= 30'b000000000000000000100110010000
                ;mem[337] <= 30'b000000000000000000100110100000
                ;mem[338] <= 30'b000000000000000000100110110000
                ;mem[339] <= 30'b000000000000000000101101000000
                ;mem[340] <= 30'b000000000000000000101101010000
                ;mem[341] <= 30'b000000000000000000101101100000
                ;mem[342] <= 30'b000000000000000000101101110000
                ;mem[343] <= 30'b000000000000000000110011110000
                ;mem[344] <= 30'b000000000000000000110100000000
                ;mem[345] <= 30'b000000000000000000110100010000
                ;mem[346] <= 30'b000000000000000000110100100000
                ;mem[347] <= 30'b000000000000000000110100110000
                ;mem[348] <= 30'b000000000000000000110101000000
                ;mem[349] <= 30'b000000000000000000111010100000
                ;mem[350] <= 30'b000000000000000000111010110000
                ;mem[351] <= 30'b000000000000000000111011000000
                ;mem[352] <= 30'b000000000000000000111011010000
                ;mem[353] <= 30'b000000000000000000111011100000
                ;mem[354] <= 30'b000000000000000000111011110000
                ;mem[355] <= 30'b000000000000000000111100000000
                ;mem[356] <= 30'b000000000000000000111100010000
                ;mem[357] <= 30'b000000000000000000111100100000
                ;mem[358] <= 30'b000000001000000000000001000000
                ;mem[359] <= 30'b000000001000000000000001010000
                ;mem[360] <= 30'b000000001000000000000001100000
                ;mem[361] <= 30'b000000001000000000000001110000
                ;mem[362] <= 30'b000000001000000000000111110000
                ;mem[363] <= 30'b000000001000000000001000000000
                ;mem[364] <= 30'b000000001000000000001000010000
                ;mem[365] <= 30'b000000001000000000001000100000
                ;mem[366] <= 30'b000000001000000000001000110000
                ;mem[367] <= 30'b000000001000000000001001000000
                ;mem[368] <= 30'b000000001000000000001110100000
                ;mem[369] <= 30'b000000001000000000001110110000
                ;mem[370] <= 30'b000000001000000000001111000000
                ;mem[371] <= 30'b000000001000000000001111010000
                ;mem[372] <= 30'b000000001000000000001111100000
                ;mem[373] <= 30'b000000001000000000001111110000
                ;mem[374] <= 30'b000000001000000000010000000000
                ;mem[375] <= 30'b000000001000000000010000010000
                ;mem[376] <= 30'b000000001000000000010000100000
                ;mem[377] <= 30'b000000001000000000010101010000
                ;mem[378] <= 30'b000000001000000000010101100000
                ;mem[379] <= 30'b000000001000000000010101110000
                ;mem[380] <= 30'b000000001000000000010110000000
                ;mem[381] <= 30'b000000001000000000010110010000
                ;mem[382] <= 30'b000000001000000000010110100000
                ;mem[383] <= 30'b000000001000000000010110110000
                ;mem[384] <= 30'b000000001000000000010111000000
                ;mem[385] <= 30'b000000001000000000010111010000
                ;mem[386] <= 30'b000000001000000000010111100000
                ;mem[387] <= 30'b000000001000000000010111110000
                ;mem[388] <= 30'b000000001000000000011100010000
                ;mem[389] <= 30'b000000001000000000011100100000
                ;mem[390] <= 30'b000000001000000000011100110000
                ;mem[391] <= 30'b000000001000000000011101000000
                ;mem[392] <= 30'b000000001000000000011101010000
                ;mem[393] <= 30'b000000001000000000011101100000
                ;mem[394] <= 30'b000000001000000000011110010000
                ;mem[395] <= 30'b000000001000000000011110100000
                ;mem[396] <= 30'b000000001000000000011110110000
                ;mem[397] <= 30'b000000001000000000100011000000
                ;mem[398] <= 30'b000000001000000000100011010000
                ;mem[399] <= 30'b000000001000000000100011100000
                ;mem[400] <= 30'b000000001000000000100011110000
                ;mem[401] <= 30'b000000001000000000100100000000
                ;mem[402] <= 30'b000000001000000000100100010000
                ;mem[403] <= 30'b000000001000000000100101100000
                ;mem[404] <= 30'b000000001000000000100101110000
                ;mem[405] <= 30'b000000001000000000100110000000
                ;mem[406] <= 30'b000000001000000000101010000000
                ;mem[407] <= 30'b000000001000000000101010010000
                ;mem[408] <= 30'b000000001000000000101010100000
                ;mem[409] <= 30'b000000001000000000101010110000
                ;mem[410] <= 30'b000000001000000000101100110000
                ;mem[411] <= 30'b000000001000000000101101000000
                ;mem[412] <= 30'b000000001000000000101101010000
                ;mem[413] <= 30'b000000001000000000110001000000
                ;mem[414] <= 30'b000000001000000000110001010000
                ;mem[415] <= 30'b000000001000000000110001100000
                ;mem[416] <= 30'b000000001000000000110011110000
                ;mem[417] <= 30'b000000001000000000110100000000
                ;mem[418] <= 30'b000000001000000000110100010000
                ;mem[419] <= 30'b000000001000000000111000000000
                ;mem[420] <= 30'b000000001000000000111000010000
                ;mem[421] <= 30'b000000001000000000111010110000
                ;mem[422] <= 30'b000000001000000000111011000000
                ;mem[423] <= 30'b000000001000000000111011010000
                ;mem[424] <= 30'b000000001000000000111011100000
                ;mem[425] <= 30'b000000001000000000111110110000
                ;mem[426] <= 30'b000000001000000000111111000000
                ;mem[427] <= 30'b000000001000000000111111010000
                ;mem[428] <= 30'b000000010000000000000000110000
                ;mem[429] <= 30'b000000010000000000000001000000
                ;mem[430] <= 30'b000000010000000000000001010000
                ;mem[431] <= 30'b000000010000000000000101000000
                ;mem[432] <= 30'b000000010000000000000101010000
                ;mem[433] <= 30'b000000010000000000000101100000
                ;mem[434] <= 30'b000000010000000000000111110000
                ;mem[435] <= 30'b000000010000000000001000000000
                ;mem[436] <= 30'b000000010000000000001000010000
                ;mem[437] <= 30'b000000010000000000001100000000
                ;mem[438] <= 30'b000000010000000000001100010000
                ;mem[439] <= 30'b000000010000000000001110110000
                ;mem[440] <= 30'b000000010000000000001111000000
                ;mem[441] <= 30'b000000010000000000001111010000
                ;mem[442] <= 30'b000000010000000000001111100000
                ;mem[443] <= 30'b000000010000000000010010110000
                ;mem[444] <= 30'b000000010000000000010011000000
                ;mem[445] <= 30'b000000010000000000010011010000
                ;mem[446] <= 30'b000000010000000000010101110000
                ;mem[447] <= 30'b000000010000000000010110000000
                ;mem[448] <= 30'b000000010000000000010110010000
                ;mem[449] <= 30'b000000010000000000011001110000
                ;mem[450] <= 30'b000000010000000000011010000000
                ;mem[451] <= 30'b000000010000000000011010010000
                ;mem[452] <= 30'b000000010000000000011100100000
                ;mem[453] <= 30'b000000010000000000011100110000
                ;mem[454] <= 30'b000000010000000000011101000000
                ;mem[455] <= 30'b000000010000000000011101010000
                ;mem[456] <= 30'b000000010000000000100000110000
                ;mem[457] <= 30'b000000010000000000100001000000
                ;mem[458] <= 30'b000000010000000000100001010000
                ;mem[459] <= 30'b000000010000000000100011000000
                ;mem[460] <= 30'b000000010000000000100011010000
                ;mem[461] <= 30'b000000010000000000100011100000
                ;mem[462] <= 30'b000000010000000000100011110000
                ;mem[463] <= 30'b000000010000000000100100000000
                ;mem[464] <= 30'b000000010000000000100111110000
                ;mem[465] <= 30'b000000010000000000101000000000
                ;mem[466] <= 30'b000000010000000000101000010000
                ;mem[467] <= 30'b000000010000000000101001110000
                ;mem[468] <= 30'b000000010000000000101010000000
                ;mem[469] <= 30'b000000010000000000101010010000
                ;mem[470] <= 30'b000000010000000000101010100000
                ;mem[471] <= 30'b000000010000000000101010110000
                ;mem[472] <= 30'b000000010000000000101011000000
                ;mem[473] <= 30'b000000010000000000101110110000
                ;mem[474] <= 30'b000000010000000000101111000000
                ;mem[475] <= 30'b000000010000000000101111010000
                ;mem[476] <= 30'b000000010000000000110000000000
                ;mem[477] <= 30'b000000010000000000110000010000
                ;mem[478] <= 30'b000000010000000000110000100000
                ;mem[479] <= 30'b000000010000000000110000110000
                ;mem[480] <= 30'b000000010000000000110001000000
                ;mem[481] <= 30'b000000010000000000110001010000
                ;mem[482] <= 30'b000000010000000000110001100000
                ;mem[483] <= 30'b000000010000000000110001110000
                ;mem[484] <= 30'b000000010000000000110110000000
                ;mem[485] <= 30'b000000010000000000110110010000
                ;mem[486] <= 30'b000000010000000000110110100000
                ;mem[487] <= 30'b000000010000000000110110110000
                ;mem[488] <= 30'b000000010000000000110111000000
                ;mem[489] <= 30'b000000010000000000110111010000
                ;mem[490] <= 30'b000000010000000000110111100000
                ;mem[491] <= 30'b000000010000000000110111110000
                ;mem[492] <= 30'b000000010000000000111000000000
                ;mem[493] <= 30'b000000010000000000111000010000
                ;mem[494] <= 30'b000000010000000000111000100000
                ;mem[495] <= 30'b000000010000000000111000110000
                ;mem[496] <= 30'b000000010000000000111101000000
                ;mem[497] <= 30'b000000010000000000111101010000
                ;mem[498] <= 30'b000000010000000000111101100000
                ;mem[499] <= 30'b000000010000000000111101110000
                ;mem[500] <= 30'b000000010000000000111110000000
                ;mem[501] <= 30'b000000010000000000111110010000
                ;mem[502] <= 30'b000000010000000000111110100000
                ;mem[503] <= 30'b000000010000000000111110110000
                ;mem[504] <= 30'b000000010000000000111111000000
                ;mem[505] <= 30'b000000010000000000111111010000
                ;mem[506] <= 30'b000000000000000001000010110000
                ;mem[507] <= 30'b000000000000000001000011000000
                ;mem[508] <= 30'b000000000000000001000011010000
                ;mem[509] <= 30'b000000000000000001000100000000
                ;mem[510] <= 30'b000000000000000001000100010000
                ;mem[511] <= 30'b000000000000000001000100100000
                ;mem[512] <= 30'b000000000000000001000100110000
                ;mem[513] <= 30'b000000000000000001000101000000
                ;mem[514] <= 30'b000000000000000001000101010000
                ;mem[515] <= 30'b000000000000000001000101100000
                ;mem[516] <= 30'b000000000000000001000101110000
                ;mem[517] <= 30'b000000000000000001001010000000
                ;mem[518] <= 30'b000000000000000001001010010000
                ;mem[519] <= 30'b000000000000000001001010100000
                ;mem[520] <= 30'b000000000000000001001010110000
                ;mem[521] <= 30'b000000000000000001001011000000
                ;mem[522] <= 30'b000000000000000001001011010000
                ;mem[523] <= 30'b000000000000000001001011100000
                ;mem[524] <= 30'b000000000000000001001011110000
                ;mem[525] <= 30'b000000000000000001001100000000
                ;mem[526] <= 30'b000000000000000001001100010000
                ;mem[527] <= 30'b000000000000000001001100100000
                ;mem[528] <= 30'b000000000000000001001100110000
                ;mem[529] <= 30'b000000000000000001010001000000
                ;mem[530] <= 30'b000000000000000001010001010000
                ;mem[531] <= 30'b000000000000000001010001100000
                ;mem[532] <= 30'b000000000000000001010001110000
                ;mem[533] <= 30'b000000000000000001010010000000
                ;mem[534] <= 30'b000000000000000001010010010000
                ;mem[535] <= 30'b000000000000000001010010100000
                ;mem[536] <= 30'b000000000000000001010010110000
                ;mem[537] <= 30'b000000000000000001010011000000
                ;mem[538] <= 30'b000000000000000001010011010000
                ;mem[539] <= 30'b000000000000000001011000010000
                ;mem[540] <= 30'b000000000000000001011000100000
                ;mem[541] <= 30'b000000000000000001011000110000
                ;mem[542] <= 30'b000000000000000001011001000000
                ;mem[543] <= 30'b000000000000000001011001010000
                ;mem[544] <= 30'b000000000000000001011001100000
                ;mem[545] <= 30'b000000000000000001011001110000
                ;mem[546] <= 30'b000000000000000001011111110000
                ;mem[547] <= 30'b000000000000000001100000000000
                ;mem[548] <= 30'b000000000000000001100000010000
                ;mem[549] <= 30'b000000000000000000100101110000
                ;mem[550] <= 30'b000000000000000000101100110000
                ;mem[551] <= 30'b000000000000000000101110110000
                ;mem[552] <= 30'b000000000000000000101111000000
                ;mem[553] <= 30'b000000000000000000110011100000
                ;mem[554] <= 30'b000000000000000000110011110000
                ;mem[555] <= 30'b000000000000000000110110000000
                ;mem[556] <= 30'b000000000000000000111010100000
                ;mem[557] <= 30'b000000000000000000111010110000
                ;mem[558] <= 30'b000000000000000000111101000000
                ;mem[559] <= 30'b000000001000000000000000110000
                ;mem[560] <= 30'b000000001000000000000010110000
                ;mem[561] <= 30'b000000001000000000000011000000
                ;mem[562] <= 30'b000000001000000000000111100000
                ;mem[563] <= 30'b000000001000000000000111110000
                ;mem[564] <= 30'b000000001000000000001010000000
                ;mem[565] <= 30'b000000001000000000001110100000
                ;mem[566] <= 30'b000000001000000000001110110000
                ;mem[567] <= 30'b000000001000000000010001000000
                ;mem[568] <= 30'b000000001000000000010101010000
                ;mem[569] <= 30'b000000001000000000010101100000
                ;mem[570] <= 30'b000000001000000000010111110000
                ;mem[571] <= 30'b000000001000000000011000000000
                ;mem[572] <= 30'b000000001000000000011100000000
                ;mem[573] <= 30'b000000001000000000011100010000
                ;mem[574] <= 30'b000000001000000000011110110000
                ;mem[575] <= 30'b000000001000000000011111000000
                ;mem[576] <= 30'b000000001000000000100011000000
                ;mem[577] <= 30'b000000001000000000100011010000
                ;mem[578] <= 30'b000000001000000000100101100000
                ;mem[579] <= 30'b000000001000000000100101110000
                ;mem[580] <= 30'b000000001000000000100110000000
                ;mem[581] <= 30'b000000001000000000101001110000
                ;mem[582] <= 30'b000000001000000000101010000000
                ;mem[583] <= 30'b000000001000000000101100100000
                ;mem[584] <= 30'b000000001000000000101100110000
                ;mem[585] <= 30'b000000001000000000110000110000
                ;mem[586] <= 30'b000000001000000000110001000000
                ;mem[587] <= 30'b000000001000000000110011010000
                ;mem[588] <= 30'b000000001000000000110011100000
                ;mem[589] <= 30'b000000001000000000110011110000
                ;mem[590] <= 30'b000000001000000000110111110000
                ;mem[591] <= 30'b000000001000000000111000000000
                ;mem[592] <= 30'b000000001000000000111010010000
                ;mem[593] <= 30'b000000001000000000111010100000
                ;mem[594] <= 30'b000000001000000000111010110000
                ;mem[595] <= 30'b000000001000000000111110110000
                ;mem[596] <= 30'b000000001000000000111111000000
                ;mem[597] <= 30'b000000010000000000000000100000
                ;mem[598] <= 30'b000000010000000000000000110000
                ;mem[599] <= 30'b000000010000000000000100110000
                ;mem[600] <= 30'b000000010000000000000101000000
                ;mem[601] <= 30'b000000010000000000000111010000
                ;mem[602] <= 30'b000000010000000000000111100000
                ;mem[603] <= 30'b000000010000000000000111110000
                ;mem[604] <= 30'b000000010000000000001011110000
                ;mem[605] <= 30'b000000010000000000001100000000
                ;mem[606] <= 30'b000000010000000000001110010000
                ;mem[607] <= 30'b000000010000000000001110100000
                ;mem[608] <= 30'b000000010000000000001110110000
                ;mem[609] <= 30'b000000010000000000010010110000
                ;mem[610] <= 30'b000000010000000000010011000000
                ;mem[611] <= 30'b000000010000000000010101010000
                ;mem[612] <= 30'b000000010000000000010101100000
                ;mem[613] <= 30'b000000010000000000011001110000
                ;mem[614] <= 30'b000000010000000000011010000000
                ;mem[615] <= 30'b000000010000000000011010010000
                ;mem[616] <= 30'b000000010000000000011011100000
                ;mem[617] <= 30'b000000010000000000011011110000
                ;mem[618] <= 30'b000000010000000000011100000000
                ;mem[619] <= 30'b000000010000000000011100010000
                ;mem[620] <= 30'b000000010000000000011100100000
                ;mem[621] <= 30'b000000010000000000100001000000
                ;mem[622] <= 30'b000000010000000000100001010000
                ;mem[623] <= 30'b000000010000000000100001100000
                ;mem[624] <= 30'b000000010000000000100001110000
                ;mem[625] <= 30'b000000010000000000100010000000
                ;mem[626] <= 30'b000000010000000000100010010000
                ;mem[627] <= 30'b000000010000000000100010100000
                ;mem[628] <= 30'b000000010000000000100010110000
                ;mem[629] <= 30'b000000010000000000100011000000
                ;mem[630] <= 30'b000000010000000000100011010000
                ;mem[631] <= 30'b000000010000000000100011100000
                ;mem[632] <= 30'b000000010000000000101010000000
                ;mem[633] <= 30'b000000010000000000101010010000
                ;mem[634] <= 30'b000000010000000000101010100000
                ;mem[635] <= 30'b000000010000000000110001010000
                ;mem[636] <= 30'b000000010000000000110001100000
                ;mem[637] <= 30'b000000010000000000111000000000
                ;mem[638] <= 30'b000000010000000000111000010000
                ;mem[639] <= 30'b000000010000000000111000100000
                ;mem[640] <= 30'b000000010000000000111111010000
                ;mem[641] <= 30'b000000010000000000111111100000
                ;mem[642] <= 30'b000000000000000001000101010000
                ;mem[643] <= 30'b000000000000000001000101100000
                ;mem[644] <= 30'b000000000000000001001100000000
                ;mem[645] <= 30'b000000000000000001001100010000
                ;mem[646] <= 30'b000000000000000001001100100000
                ;mem[647] <= 30'b000000000000000001010011010000
                ;mem[648] <= 30'b000000000000000001010011100000
                ;mem[649] <= 30'b000000000000000001011010000000
                ;mem[650] <= 30'b000000000000000001011010010000
                ;mem[651] <= 30'b000000000000000001011010100000
                ;mem[652] <= 30'b000000000000000001100001000000
                ;mem[653] <= 30'b000000000000000001100001010000
                ;mem[654] <= 30'b000000000000000001101000000000
                ;mem[655] <= 30'b000000000000000000100111010000
                ;mem[656] <= 30'b000000000000000000101110000000
                ;mem[657] <= 30'b000000000000000000101110010000
                ;mem[658] <= 30'b000000000000000000101110100000
                ;mem[659] <= 30'b000000000000000000110101000000
                ;mem[660] <= 30'b000000000000000000110101010000
                ;mem[661] <= 30'b000000000000000000110101100000
                ;mem[662] <= 30'b000000000000000000111011110000
                ;mem[663] <= 30'b000000000000000000111100000000
                ;mem[664] <= 30'b000000000000000000111100010000
                ;mem[665] <= 30'b000000001000000000000010000000
                ;mem[666] <= 30'b000000001000000000000010010000
                ;mem[667] <= 30'b000000001000000000000010100000
                ;mem[668] <= 30'b000000001000000000001001000000
                ;mem[669] <= 30'b000000001000000000001001010000
                ;mem[670] <= 30'b000000001000000000001001100000
                ;mem[671] <= 30'b000000001000000000001111110000
                ;mem[672] <= 30'b000000001000000000010000000000
                ;mem[673] <= 30'b000000001000000000010000010000
                ;mem[674] <= 30'b000000001000000000010110110000
                ;mem[675] <= 30'b000000001000000000010111000000
                ;mem[676] <= 30'b000000001000000000010111010000
                ;mem[677] <= 30'b000000001000000000011101100000
                ;mem[678] <= 30'b000000001000000000011101110000
                ;mem[679] <= 30'b000000001000000000011110000000
                ;mem[680] <= 30'b000000001000000000011110010000
                ;mem[681] <= 30'b000000001000000000100100100000
                ;mem[682] <= 30'b000000001000000000100100110000
                ;mem[683] <= 30'b000000001000000000100101000000
                ;mem[684] <= 30'b000000001000000000101011100000
                ;mem[685] <= 30'b000000001000000000101011110000
                ;mem[686] <= 30'b000000001000000000101100000000
                ;mem[687] <= 30'b000000001000000000110010100000
                ;mem[688] <= 30'b000000001000000000110010110000
                ;mem[689] <= 30'b000000001000000000110011000000
                ;mem[690] <= 30'b000000001000000000111001010000
                ;mem[691] <= 30'b000000001000000000111001100000
                ;mem[692] <= 30'b000000001000000000111001110000
                ;mem[693] <= 30'b000000010000000000000000000000
                ;mem[694] <= 30'b000000010000000000000110100000
                ;mem[695] <= 30'b000000010000000000000110110000
                ;mem[696] <= 30'b000000010000000000000111000000
                ;mem[697] <= 30'b000000010000000000001101010000
                ;mem[698] <= 30'b000000010000000000001101100000
                ;mem[699] <= 30'b000000010000000000001101110000
                ;mem[700] <= 30'b000000010000000000010100010000
                ;mem[701] <= 30'b000000010000000000010100100000
                ;mem[702] <= 30'b000000010000000000010100110000
                ;mem[703] <= 30'b000000010000000000011011010000
                ;mem[704] <= 30'b000000010000000000011011100000
                ;mem[705] <= 30'b000000010000000000011011110000
                ;mem[706] <= 30'b000000010000000000100010000000
                ;mem[707] <= 30'b000000010000000000100010010000
                ;mem[708] <= 30'b000000010000000000100010100000
                ;mem[709] <= 30'b000000010000000000101001000000
                ;mem[710] <= 30'b000000010000000000101001010000
                ;mem[711] <= 30'b000000010000000000101001100000
                ;mem[712] <= 30'b000000010000000000110000000000
                ;mem[713] <= 30'b000000010000000000110000010000
                ;mem[714] <= 30'b000000010000000000110000100000
                ;mem[715] <= 30'b000000010000000000110111000000
                ;mem[716] <= 30'b000000010000000000110111010000
                ;mem[717] <= 30'b000000010000000000111101110000
                ;mem[718] <= 30'b000000010000000000111110000000
                ;mem[719] <= 30'b000000010000000000111110010000
                ;mem[720] <= 30'b000000000000000001000100000000
                ;mem[721] <= 30'b000000000000000001000100010000
                ;mem[722] <= 30'b000000000000000001000100100000
                ;mem[723] <= 30'b000000000000000001001011000000
                ;mem[724] <= 30'b000000000000000001001011010000
                ;mem[725] <= 30'b000000000000000001010001110000
                ;mem[726] <= 30'b000000000000000001010010000000
                ;mem[727] <= 30'b000000000000000001010010010000
                ;mem[728] <= 30'b000000000000000001011000110000
                ;mem[729] <= 30'b000000000000000001011001000000
                ;mem[730] <= 30'b000000000000000001011001010000
                ;mem[731] <= 30'b000000000000000001011111110000
                ;mem[732] <= 30'b000000000000000001100000000000
                ;mem[733] <= 30'b000000000000000001100000010000
                ;mem[734] <= 30'b000000000000000001100111000000
                ;mem[735] <= 30'b000000000000000000100101100000
                ;mem[736] <= 30'b000000000000000000100101110000
                ;mem[737] <= 30'b000000000000000000101100010000
                ;mem[738] <= 30'b000000000000000000101100100000
                ;mem[739] <= 30'b000000000000000000101100110000
                ;mem[740] <= 30'b000000000000000000101111010000
                ;mem[741] <= 30'b000000000000000000101111100000
                ;mem[742] <= 30'b000000000000000000110011000000
                ;mem[743] <= 30'b000000000000000000110011010000
                ;mem[744] <= 30'b000000000000000000110011100000
                ;mem[745] <= 30'b000000000000000000110110000000
                ;mem[746] <= 30'b000000000000000000110110010000
                ;mem[747] <= 30'b000000000000000000111010000000
                ;mem[748] <= 30'b000000000000000000111010010000
                ;mem[749] <= 30'b000000000000000000111101000000
                ;mem[750] <= 30'b000000000000000000111101010000
                ;mem[751] <= 30'b000000001000000000000000010000
                ;mem[752] <= 30'b000000001000000000000000100000
                ;mem[753] <= 30'b000000001000000000000000110000
                ;mem[754] <= 30'b000000001000000000000011010000
                ;mem[755] <= 30'b000000001000000000000011100000
                ;mem[756] <= 30'b000000001000000000000111000000
                ;mem[757] <= 30'b000000001000000000000111010000
                ;mem[758] <= 30'b000000001000000000000111100000
                ;mem[759] <= 30'b000000001000000000001010000000
                ;mem[760] <= 30'b000000001000000000001010010000
                ;mem[761] <= 30'b000000001000000000001110000000
                ;mem[762] <= 30'b000000001000000000001110010000
                ;mem[763] <= 30'b000000001000000000010001000000
                ;mem[764] <= 30'b000000001000000000010001010000
                ;mem[765] <= 30'b000000001000000000010100110000
                ;mem[766] <= 30'b000000001000000000010101000000
                ;mem[767] <= 30'b000000001000000000010111110000
                ;mem[768] <= 30'b000000001000000000011000000000
                ;mem[769] <= 30'b000000001000000000011011100000
                ;mem[770] <= 30'b000000001000000000011011110000
                ;mem[771] <= 30'b000000001000000000011100000000
                ;mem[772] <= 30'b000000001000000000011110110000
                ;mem[773] <= 30'b000000001000000000011111000000
                ;mem[774] <= 30'b000000001000000000100010100000
                ;mem[775] <= 30'b000000001000000000100010110000
                ;mem[776] <= 30'b000000001000000000100011000000
                ;mem[777] <= 30'b000000001000000000100101010000
                ;mem[778] <= 30'b000000001000000000100101100000
                ;mem[779] <= 30'b000000001000000000100101110000
                ;mem[780] <= 30'b000000001000000000101001100000
                ;mem[781] <= 30'b000000001000000000101001110000
                ;mem[782] <= 30'b000000001000000000101010000000
                ;mem[783] <= 30'b000000001000000000101010010000
                ;mem[784] <= 30'b000000001000000000101010100000
                ;mem[785] <= 30'b000000001000000000101011110000
                ;mem[786] <= 30'b000000001000000000101100000000
                ;mem[787] <= 30'b000000001000000000101100010000
                ;mem[788] <= 30'b000000001000000000101100100000
                ;mem[789] <= 30'b000000001000000000101100110000
                ;mem[790] <= 30'b000000001000000000110000110000
                ;mem[791] <= 30'b000000001000000000110001000000
                ;mem[792] <= 30'b000000001000000000110001010000
                ;mem[793] <= 30'b000000001000000000110001100000
                ;mem[794] <= 30'b000000001000000000110001110000
                ;mem[795] <= 30'b000000001000000000110010000000
                ;mem[796] <= 30'b000000001000000000110010010000
                ;mem[797] <= 30'b000000001000000000110010100000
                ;mem[798] <= 30'b000000001000000000110010110000
                ;mem[799] <= 30'b000000001000000000110011000000
                ;mem[800] <= 30'b000000001000000000110011010000
                ;mem[801] <= 30'b000000001000000000110011100000
                ;mem[802] <= 30'b000000001000000000111000010000
                ;mem[803] <= 30'b000000001000000000111000100000
                ;mem[804] <= 30'b000000001000000000111000110000
                ;mem[805] <= 30'b000000001000000000111001000000
                ;mem[806] <= 30'b000000001000000000111001010000
                ;mem[807] <= 30'b000000001000000000111001100000
                ;mem[808] <= 30'b000000001000000000111010000000
                ;mem[809] <= 30'b000000001000000000111010010000
                ;mem[810] <= 30'b000000001000000000111010100000
                ;mem[811] <= 30'b000000010000000000000000000000
                ;mem[812] <= 30'b000000010000000000000000010000
                ;mem[813] <= 30'b000000010000000000000000100000
                ;mem[814] <= 30'b000000010000000000000000110000
                ;mem[815] <= 30'b000000010000000000000100110000
                ;mem[816] <= 30'b000000010000000000000101000000
                ;mem[817] <= 30'b000000010000000000000101010000
                ;mem[818] <= 30'b000000010000000000000101100000
                ;mem[819] <= 30'b000000010000000000000101110000
                ;mem[820] <= 30'b000000010000000000000110000000
                ;mem[821] <= 30'b000000010000000000000110010000
                ;mem[822] <= 30'b000000010000000000000110100000
                ;mem[823] <= 30'b000000010000000000000110110000
                ;mem[824] <= 30'b000000010000000000000111000000
                ;mem[825] <= 30'b000000010000000000000111010000
                ;mem[826] <= 30'b000000010000000000000111100000
                ;mem[827] <= 30'b000000010000000000001100010000
                ;mem[828] <= 30'b000000010000000000001100100000
                ;mem[829] <= 30'b000000010000000000001100110000
                ;mem[830] <= 30'b000000010000000000001101000000
                ;mem[831] <= 30'b000000010000000000001101010000
                ;mem[832] <= 30'b000000010000000000001101100000
                ;mem[833] <= 30'b000000010000000000001110000000
                ;mem[834] <= 30'b000000010000000000001110010000
                ;mem[835] <= 30'b000000010000000000001110100000
                ;mem[836] <= 30'b000000010000000000010101000000
                ;mem[837] <= 30'b000000010000000000010101010000
                ;mem[838] <= 30'b000000010000000000011011110000
                ;mem[839] <= 30'b000000010000000000011100000000
                ;mem[840] <= 30'b000000010000000000100010110000
                ;mem[841] <= 30'b000000010000000000100011000000
                ;mem[842] <= 30'b000000010000000000101001100000
                ;mem[843] <= 30'b000000010000000000101001110000
                ;mem[844] <= 30'b000000010000000000101010000000
                ;mem[845] <= 30'b000000010000000000110000100000
                ;mem[846] <= 30'b000000010000000000110000110000
                ;mem[847] <= 30'b000000010000000000110111100000
                ;mem[848] <= 30'b000000010000000000110111110000
                ;mem[849] <= 30'b000000010000000000111110010000
                ;mem[850] <= 30'b000000010000000000111110100000
                ;mem[851] <= 30'b000000010000000000111110110000
                ;mem[852] <= 30'b000000000000000001000100100000
                ;mem[853] <= 30'b000000000000000001000100110000
                ;mem[854] <= 30'b000000000000000001001011100000
                ;mem[855] <= 30'b000000000000000001001011110000
                ;mem[856] <= 30'b000000000000000001010010010000
                ;mem[857] <= 30'b000000000000000001010010100000
                ;mem[858] <= 30'b000000000000000001010010110000
                ;mem[859] <= 30'b000000000000000001011001010000
                ;mem[860] <= 30'b000000000000000001011001100000
                ;mem[861] <= 30'b000000000000000001011001110000
                ;mem[862] <= 30'b000000000000000001011010010000
                ;mem[863] <= 30'b000000000000000001011010100000
                ;mem[864] <= 30'b000000000000000001100000010000
                ;mem[865] <= 30'b000000000000000001100000100000
                ;mem[866] <= 30'b000000000000000001100000110000
                ;mem[867] <= 30'b000000000000000001100001000000
                ;mem[868] <= 30'b000000000000000001100001010000
                ;mem[869] <= 30'b000000000000000001100111100000
                ;mem[870] <= 30'b000000000000000001100111110000
                ;mem[871] <= 30'b000000000000000000101101000000
                ;mem[872] <= 30'b000000000000000000101101010000
                ;mem[873] <= 30'b000000000000000000110011110000
                ;mem[874] <= 30'b000000000000000000110100000000
                ;mem[875] <= 30'b000000000000000000110100010000
                ;mem[876] <= 30'b000000000000000000111010100000
                ;mem[877] <= 30'b000000000000000000111010110000
                ;mem[878] <= 30'b000000000000000000111011000000
                ;mem[879] <= 30'b000000000000000000111011010000
                ;mem[880] <= 30'b000000000000000000111011100000
                ;mem[881] <= 30'b000000001000000000000001000000
                ;mem[882] <= 30'b000000001000000000000001010000
                ;mem[883] <= 30'b000000001000000000000111110000
                ;mem[884] <= 30'b000000001000000000001000000000
                ;mem[885] <= 30'b000000001000000000001000010000
                ;mem[886] <= 30'b000000001000000000001110100000
                ;mem[887] <= 30'b000000001000000000001110110000
                ;mem[888] <= 30'b000000001000000000001111000000
                ;mem[889] <= 30'b000000001000000000001111010000
                ;mem[890] <= 30'b000000001000000000001111100000
                ;mem[891] <= 30'b000000001000000000010101010000
                ;mem[892] <= 30'b000000001000000000010101100000
                ;mem[893] <= 30'b000000001000000000010101110000
                ;mem[894] <= 30'b000000001000000000010110000000
                ;mem[895] <= 30'b000000001000000000010110010000
                ;mem[896] <= 30'b000000001000000000010110100000
                ;mem[897] <= 30'b000000001000000000010110110000
                ;mem[898] <= 30'b000000001000000000011100010000
                ;mem[899] <= 30'b000000001000000000011100100000
                ;mem[900] <= 30'b000000001000000000011100110000
                ;mem[901] <= 30'b000000001000000000011101000000
                ;mem[902] <= 30'b000000001000000000011101010000
                ;mem[903] <= 30'b000000001000000000011101100000
                ;mem[904] <= 30'b000000001000000000011101110000
                ;mem[905] <= 30'b000000001000000000011110000000
                ;mem[906] <= 30'b000000001000000000100011010000
                ;mem[907] <= 30'b000000001000000000100011100000
                ;mem[908] <= 30'b000000001000000000100100100000
                ;mem[909] <= 30'b000000001000000000100100110000
                ;mem[910] <= 30'b000000001000000000100101000000
                ;mem[911] <= 30'b000000001000000000100101010000
                ;mem[912] <= 30'b000000001000000000101010010000
                ;mem[913] <= 30'b000000001000000000101011100000
                ;mem[914] <= 30'b000000001000000000101011110000
                ;mem[915] <= 30'b000000001000000000101100000000
                ;mem[916] <= 30'b000000001000000000101100010000
                ;mem[917] <= 30'b000000001000000000110001000000
                ;mem[918] <= 30'b000000001000000000110001010000
                ;mem[919] <= 30'b000000001000000000110001100000
                ;mem[920] <= 30'b000000001000000000110010100000
                ;mem[921] <= 30'b000000001000000000110010110000
                ;mem[922] <= 30'b000000001000000000110011000000
                ;mem[923] <= 30'b000000001000000000110011010000
                ;mem[924] <= 30'b000000001000000000111000010000
                ;mem[925] <= 30'b000000001000000000111000100000
                ;mem[926] <= 30'b000000001000000000111001010000
                ;mem[927] <= 30'b000000001000000000111001100000
                ;mem[928] <= 30'b000000001000000000111001110000
                ;mem[929] <= 30'b000000001000000000111010000000
                ;mem[930] <= 30'b000000001000000000111010010000
                ;mem[931] <= 30'b000000001000000000111111010000
                ;mem[932] <= 30'b000000001000000000111111100000
                ;mem[933] <= 30'b000000001000000000111111110000
                ;mem[934] <= 30'b000000010000000000000000000000
                ;mem[935] <= 30'b000000010000000000000000010000
                ;mem[936] <= 30'b000000010000000000000101000000
                ;mem[937] <= 30'b000000010000000000000101010000
                ;mem[938] <= 30'b000000010000000000000101100000
                ;mem[939] <= 30'b000000010000000000000110100000
                ;mem[940] <= 30'b000000010000000000000110110000
                ;mem[941] <= 30'b000000010000000000000111000000
                ;mem[942] <= 30'b000000010000000000000111010000
                ;mem[943] <= 30'b000000010000000000001100010000
                ;mem[944] <= 30'b000000010000000000001100100000
                ;mem[945] <= 30'b000000010000000000001101010000
                ;mem[946] <= 30'b000000010000000000001101100000
                ;mem[947] <= 30'b000000010000000000001101110000
                ;mem[948] <= 30'b000000010000000000001110000000
                ;mem[949] <= 30'b000000010000000000001110010000
                ;mem[950] <= 30'b000000010000000000010011010000
                ;mem[951] <= 30'b000000010000000000010011100000
                ;mem[952] <= 30'b000000010000000000010011110000
                ;mem[953] <= 30'b000000010000000000010100000000
                ;mem[954] <= 30'b000000010000000000010100010000
                ;mem[955] <= 30'b000000010000000000010100100000
                ;mem[956] <= 30'b000000010000000000010101000000
                ;mem[957] <= 30'b000000010000000000010101010000
                ;mem[958] <= 30'b000000010000000000010101100000
                ;mem[959] <= 30'b000000010000000000011010100000
                ;mem[960] <= 30'b000000010000000000011010110000
                ;mem[961] <= 30'b000000010000000000011011000000
                ;mem[962] <= 30'b000000010000000000011011010000
                ;mem[963] <= 30'b000000010000000000011100000000
                ;mem[964] <= 30'b000000010000000000011100010000
                ;mem[965] <= 30'b000000010000000000011100100000
                ;mem[966] <= 30'b000000010000000000100001110000
                ;mem[967] <= 30'b000000010000000000100010000000
                ;mem[968] <= 30'b000000010000000000100011010000
                ;mem[969] <= 30'b000000010000000000100011100000
                ;mem[970] <= 30'b000000010000000000100011110000
                ;mem[971] <= 30'b000000010000000000101010100000
                ;mem[972] <= 30'b000000010000000000101010110000
                ;mem[973] <= 30'b000000010000000000110001100000
                ;mem[974] <= 30'b000000010000000000110001110000
                ;mem[975] <= 30'b000000010000000000111000110000
                ;mem[976] <= 30'b000000010000000000111001000000
                ;mem[977] <= 30'b000000000000000001000101100000
                ;mem[978] <= 30'b000000000000000001000101110000
                ;mem[979] <= 30'b000000000000000001001100110000
                ;mem[980] <= 30'b000000000000000001001101000000
                ;mem[981] <= 30'b000000000000000001010100000000
                ;mem[982] <= 30'b000000000000000001010100010000
                ;mem[983] <= 30'b000000000000000001011011000000
                ;mem[984] <= 30'b000000000000000001011011010000
                ;mem[985] <= 30'b000000000000000001100010010000
                ;mem[986] <= 30'b000000000000000001100010100000
                ;mem[987] <= 30'b000000000000000001101001010000
                ;mem[988] <= 30'b000000000000000001101001100000
                ;mem[989] <= 30'b000000000000000001110000100000
                ;mem[990] <= 30'b000000000000000000100001100000
                ;mem[991] <= 30'b000000000000000000100111000000
                ;mem[992] <= 30'b000000000000000000100111010000
                ;mem[993] <= 30'b000000000000000000100111100000
                ;mem[994] <= 30'b000000000000000000100111110000
                ;mem[995] <= 30'b000000000000000000101000000000
                ;mem[996] <= 30'b000000000000000000101000010000
                ;mem[997] <= 30'b000000000000000000101000100000
                ;mem[998] <= 30'b000000000000000000101000110000
                ;mem[999] <= 30'b000000000000000000101001000000
                ;mem[1000] <= 30'b000000000000000000101101010000
                ;mem[1001] <= 30'b000000000000000000101101100000
                ;mem[1002] <= 30'b000000000000000000101101110000
                ;mem[1003] <= 30'b000000000000000000101110000000
                ;mem[1004] <= 30'b000000000000000000101110010000
                ;mem[1005] <= 30'b000000000000000000101110100000
                ;mem[1006] <= 30'b000000000000000000101110110000
                ;mem[1007] <= 30'b000000000000000000101111000000
                ;mem[1008] <= 30'b000000000000000000101111010000
                ;mem[1009] <= 30'b000000000000000000101111100000
                ;mem[1010] <= 30'b000000000000000000101111110000
                ;mem[1011] <= 30'b000000000000000000110000000000
                ;mem[1012] <= 30'b000000000000000000110100010000
                ;mem[1013] <= 30'b000000000000000000110100100000
                ;mem[1014] <= 30'b000000000000000000110100110000
                ;mem[1015] <= 30'b000000000000000000110101000000
                ;mem[1016] <= 30'b000000000000000000110101010000
                ;mem[1017] <= 30'b000000000000000000110101100000
                ;mem[1018] <= 30'b000000000000000000110101110000
                ;mem[1019] <= 30'b000000000000000000110110000000
                ;mem[1020] <= 30'b000000000000000000110110010000
                ;mem[1021] <= 30'b000000000000000000110110100000
                ;mem[1022] <= 30'b000000000000000000110110110000
                ;mem[1023] <= 30'b000000000000000000110111000000
                ;mem[1024] <= 30'b000000000000000000111010010000
                ;mem[1025] <= 30'b000000000000000000111011010000
                ;mem[1026] <= 30'b000000000000000000111011100000
                ;mem[1027] <= 30'b000000000000000000111011110000
                ;mem[1028] <= 30'b000000000000000000111100000000
                ;mem[1029] <= 30'b000000001000000000000001010000
                ;mem[1030] <= 30'b000000001000000000000001100000
                ;mem[1031] <= 30'b000000001000000000000001110000
                ;mem[1032] <= 30'b000000001000000000000010000000
                ;mem[1033] <= 30'b000000001000000000000010010000
                ;mem[1034] <= 30'b000000001000000000000010100000
                ;mem[1035] <= 30'b000000001000000000000010110000
                ;mem[1036] <= 30'b000000001000000000000011000000
                ;mem[1037] <= 30'b000000001000000000000011010000
                ;mem[1038] <= 30'b000000001000000000000011100000
                ;mem[1039] <= 30'b000000001000000000000011110000
                ;mem[1040] <= 30'b000000001000000000000100000000
                ;mem[1041] <= 30'b000000001000000000001000010000
                ;mem[1042] <= 30'b000000001000000000001000100000
                ;mem[1043] <= 30'b000000001000000000001000110000
                ;mem[1044] <= 30'b000000001000000000001001000000
                ;mem[1045] <= 30'b000000001000000000001001010000
                ;mem[1046] <= 30'b000000001000000000001001100000
                ;mem[1047] <= 30'b000000001000000000001001110000
                ;mem[1048] <= 30'b000000001000000000001010000000
                ;mem[1049] <= 30'b000000001000000000001010010000
                ;mem[1050] <= 30'b000000001000000000001010100000
                ;mem[1051] <= 30'b000000001000000000001010110000
                ;mem[1052] <= 30'b000000001000000000001011000000
                ;mem[1053] <= 30'b000000001000000000001110010000
                ;mem[1054] <= 30'b000000001000000000001111010000
                ;mem[1055] <= 30'b000000001000000000001111100000
                ;mem[1056] <= 30'b000000001000000000001111110000
                ;mem[1057] <= 30'b000000001000000000010000000000
                ;mem[1058] <= 30'b000000001000000000010101000000
                ;mem[1059] <= 30'b000000001000000000010101010000
                ;mem[1060] <= 30'b000000001000000000011011110000
                ;mem[1061] <= 30'b000000001000000000011100000000
                ;mem[1062] <= 30'b000000001000000000011100010000
                ;mem[1063] <= 30'b000000001000000000100010100000
                ;mem[1064] <= 30'b000000001000000000100010110000
                ;mem[1065] <= 30'b000000001000000000100011000000
                ;mem[1066] <= 30'b000000001000000000101001100000
                ;mem[1067] <= 30'b000000001000000000101001110000
                ;mem[1068] <= 30'b000000001000000000110000010000
                ;mem[1069] <= 30'b000000001000000000110000100000
                ;mem[1070] <= 30'b000000001000000000110000110000
                ;mem[1071] <= 30'b000000001000000000110111010000
                ;mem[1072] <= 30'b000000001000000000110111100000
                ;mem[1073] <= 30'b000000001000000000110111110000
                ;mem[1074] <= 30'b000000001000000000111110010000
                ;mem[1075] <= 30'b000000001000000000111110100000
                ;mem[1076] <= 30'b000000001000000000111110110000
                ;mem[1077] <= 30'b000000001000000000111111000000
                ;mem[1078] <= 30'b000000001000000000111111010000
                ;mem[1079] <= 30'b000000001000000000111111100000
                ;mem[1080] <= 30'b000000010000000000000100010000
                ;mem[1081] <= 30'b000000010000000000000100100000
                ;mem[1082] <= 30'b000000010000000000000100110000
                ;mem[1083] <= 30'b000000010000000000001011010000
                ;mem[1084] <= 30'b000000010000000000001011100000
                ;mem[1085] <= 30'b000000010000000000001011110000
                ;mem[1086] <= 30'b000000010000000000010010010000
                ;mem[1087] <= 30'b000000010000000000010010100000
                ;mem[1088] <= 30'b000000010000000000010010110000
                ;mem[1089] <= 30'b000000010000000000010011000000
                ;mem[1090] <= 30'b000000010000000000010011010000
                ;mem[1091] <= 30'b000000010000000000010011100000
                ;mem[1092] <= 30'b000000010000000000011001010000
                ;mem[1093] <= 30'b000000010000000000011001100000
                ;mem[1094] <= 30'b000000010000000000011001110000
                ;mem[1095] <= 30'b000000010000000000011010000000
                ;mem[1096] <= 30'b000000010000000000011010010000
                ;mem[1097] <= 30'b000000010000000000011010100000
                ;mem[1098] <= 30'b000000010000000000011010110000
                ;mem[1099] <= 30'b000000010000000000011011000000
                ;mem[1100] <= 30'b000000010000000000011011010000
                ;mem[1101] <= 30'b000000010000000000011011100000
                ;mem[1102] <= 30'b000000010000000000011011110000
                ;mem[1103] <= 30'b000000010000000000011100000000
                ;mem[1104] <= 30'b000000010000000000011100010000
                ;mem[1105] <= 30'b000000010000000000011100100000
                ;mem[1106] <= 30'b000000010000000000100000110000
                ;mem[1107] <= 30'b000000010000000000100001000000
                ;mem[1108] <= 30'b000000010000000000100001010000
                ;mem[1109] <= 30'b000000010000000000100001100000
                ;mem[1110] <= 30'b000000010000000000100001110000
                ;mem[1111] <= 30'b000000010000000000100010000000
                ;mem[1112] <= 30'b000000010000000000100010010000
                ;mem[1113] <= 30'b000000010000000000100010100000
                ;mem[1114] <= 30'b000000010000000000100010110000
                ;mem[1115] <= 30'b000000010000000000100011000000
                ;mem[1116] <= 30'b000000010000000000100011010000
                ;mem[1117] <= 30'b000000010000000000100011100000
                ;mem[1118] <= 30'b000000010000000000101000110000
                ;mem[1119] <= 30'b000000010000000000101001000000
                ;mem[1120] <= 30'b000000010000000000101001010000
                ;mem[1121] <= 30'b000000010000000000101001100000
                ;mem[1122] <= 30'b000000010000000000101001110000
                ;mem[1123] <= 30'b000000010000000000101010000000
                ;mem[1124] <= 30'b000000010000000000101010010000
                ;mem[1125] <= 30'b000000010000000000101010100000
                ;mem[1126] <= 30'b000000010000000000101010110000
                ;mem[1127] <= 30'b000000010000000000110000000000
                ;mem[1128] <= 30'b000000010000000000110000010000
                ;mem[1129] <= 30'b000000010000000000110000100000
                ;mem[1130] <= 30'b000000010000000000110001000000
                ;mem[1131] <= 30'b000000010000000000110001010000
                ;mem[1132] <= 30'b000000010000000000110001100000
                ;mem[1133] <= 30'b000000010000000000110001110000
                ;mem[1134] <= 30'b000000010000000000110111000000
                ;mem[1135] <= 30'b000000010000000000110111010000
                ;mem[1136] <= 30'b000000010000000000110111100000
                ;mem[1137] <= 30'b000000010000000000110111110000
                ;mem[1138] <= 30'b000000010000000000111000000000
                ;mem[1139] <= 30'b000000010000000000111000010000
                ;mem[1140] <= 30'b000000010000000000111000100000
                ;mem[1141] <= 30'b000000010000000000111000110000
                ;mem[1142] <= 30'b000000010000000000111110000000
                ;mem[1143] <= 30'b000000010000000000111110010000
                ;mem[1144] <= 30'b000000010000000000111110100000
                ;mem[1145] <= 30'b000000010000000000111110110000
                ;mem[1146] <= 30'b000000010000000000111111000000
                ;mem[1147] <= 30'b000000010000000000111111010000
                ;mem[1148] <= 30'b000000010000000000111111100000
                ;mem[1149] <= 30'b000000000000000001000100000000
                ;mem[1150] <= 30'b000000000000000001000100010000
                ;mem[1151] <= 30'b000000000000000001000100100000
                ;mem[1152] <= 30'b000000000000000001000101000000
                ;mem[1153] <= 30'b000000000000000001000101010000
                ;mem[1154] <= 30'b000000000000000001000101100000
                ;mem[1155] <= 30'b000000000000000001000101110000
                ;mem[1156] <= 30'b000000000000000001001011000000
                ;mem[1157] <= 30'b000000000000000001001011010000
                ;mem[1158] <= 30'b000000000000000001001011100000
                ;mem[1159] <= 30'b000000000000000001001011110000
                ;mem[1160] <= 30'b000000000000000001001100000000
                ;mem[1161] <= 30'b000000000000000001001100010000
                ;mem[1162] <= 30'b000000000000000001001100100000
                ;mem[1163] <= 30'b000000000000000001001100110000
                ;mem[1164] <= 30'b000000000000000001010010000000
                ;mem[1165] <= 30'b000000000000000001010010010000
                ;mem[1166] <= 30'b000000000000000001010010100000
                ;mem[1167] <= 30'b000000000000000001010010110000
                ;mem[1168] <= 30'b000000000000000001010011000000
                ;mem[1169] <= 30'b000000000000000001010011010000
                ;mem[1170] <= 30'b000000000000000001010011100000
                ;mem[1171] <= 30'b000000000000000001011001010000
                ;mem[1172] <= 30'b000000000000000001011001100000
                ;mem[1173] <= 30'b000000000000000001011001110000
                ;mem[1174] <= 30'b000000000000000001011010000000
                ;mem[1175] <= 30'b000000000000000001011010010000
                ;mem[1176] <= 30'b000000000000000001100000110000
                ;mem[1177] <= 30'b000000000000000000110100110000
                ;mem[1178] <= 30'b000000000000000000110101000000
                ;mem[1179] <= 30'b000000000000000000110101010000
                ;mem[1180] <= 30'b000000000000000000111011000000
                ;mem[1181] <= 30'b000000000000000000111011010000
                ;mem[1182] <= 30'b000000000000000000111011100000
                ;mem[1183] <= 30'b000000000000000000111011110000
                ;mem[1184] <= 30'b000000000000000000111100000000
                ;mem[1185] <= 30'b000000000000000000111100010000
                ;mem[1186] <= 30'b000000000000000000111100100000
                ;mem[1187] <= 30'b000000000000000000111100110000
                ;mem[1188] <= 30'b000000000000000000111101000000
                ;mem[1189] <= 30'b000000000000000000111101010000
                ;mem[1190] <= 30'b000000001000000000001000110000
                ;mem[1191] <= 30'b000000001000000000001001000000
                ;mem[1192] <= 30'b000000001000000000001001010000
                ;mem[1193] <= 30'b000000001000000000001111000000
                ;mem[1194] <= 30'b000000001000000000001111010000
                ;mem[1195] <= 30'b000000001000000000001111100000
                ;mem[1196] <= 30'b000000001000000000001111110000
                ;mem[1197] <= 30'b000000001000000000010000000000
                ;mem[1198] <= 30'b000000001000000000010000010000
                ;mem[1199] <= 30'b000000001000000000010000100000
                ;mem[1200] <= 30'b000000001000000000010000110000
                ;mem[1201] <= 30'b000000001000000000010001000000
                ;mem[1202] <= 30'b000000001000000000010001010000
                ;mem[1203] <= 30'b000000001000000000010101100000
                ;mem[1204] <= 30'b000000001000000000010101110000
                ;mem[1205] <= 30'b000000001000000000010110000000
                ;mem[1206] <= 30'b000000001000000000010110010000
                ;mem[1207] <= 30'b000000001000000000010110100000
                ;mem[1208] <= 30'b000000001000000000010110110000
                ;mem[1209] <= 30'b000000001000000000010111000000
                ;mem[1210] <= 30'b000000001000000000010111010000
                ;mem[1211] <= 30'b000000001000000000010111100000
                ;mem[1212] <= 30'b000000001000000000010111110000
                ;mem[1213] <= 30'b000000001000000000011000000000
                ;mem[1214] <= 30'b000000001000000000011000010000
                ;mem[1215] <= 30'b000000001000000000011100000000
                ;mem[1216] <= 30'b000000001000000000011100010000
                ;mem[1217] <= 30'b000000001000000000011100100000
                ;mem[1218] <= 30'b000000001000000000011100110000
                ;mem[1219] <= 30'b000000001000000000011101000000
                ;mem[1220] <= 30'b000000001000000000011101010000
                ;mem[1221] <= 30'b000000001000000000011110010000
                ;mem[1222] <= 30'b000000001000000000011110110000
                ;mem[1223] <= 30'b000000001000000000011111000000
                ;mem[1224] <= 30'b000000001000000000011111010000
                ;mem[1225] <= 30'b000000001000000000011111100000
                ;mem[1226] <= 30'b000000001000000000100011000000
                ;mem[1227] <= 30'b000000001000000000100011010000
                ;mem[1228] <= 30'b000000001000000000100011100000
                ;mem[1229] <= 30'b000000001000000000100011110000
                ;mem[1230] <= 30'b000000001000000000100101010000
                ;mem[1231] <= 30'b000000001000000000100110000000
                ;mem[1232] <= 30'b000000001000000000100110010000
                ;mem[1233] <= 30'b000000001000000000100110100000
                ;mem[1234] <= 30'b000000001000000000101001110000
                ;mem[1235] <= 30'b000000001000000000101010000000
                ;mem[1236] <= 30'b000000001000000000101010010000
                ;mem[1237] <= 30'b000000001000000000101100100000
                ;mem[1238] <= 30'b000000001000000000101100110000
                ;mem[1239] <= 30'b000000001000000000101101000000
                ;mem[1240] <= 30'b000000001000000000101101010000
                ;mem[1241] <= 30'b000000001000000000101101100000
                ;mem[1242] <= 30'b000000001000000000110000110000
                ;mem[1243] <= 30'b000000001000000000110001000000
                ;mem[1244] <= 30'b000000001000000000110001010000
                ;mem[1245] <= 30'b000000001000000000110001110000
                ;mem[1246] <= 30'b000000001000000000110010000000
                ;mem[1247] <= 30'b000000001000000000110010010000
                ;mem[1248] <= 30'b000000001000000000110010100000
                ;mem[1249] <= 30'b000000001000000000110010110000
                ;mem[1250] <= 30'b000000001000000000110011000000
                ;mem[1251] <= 30'b000000001000000000110011010000
                ;mem[1252] <= 30'b000000001000000000110011100000
                ;mem[1253] <= 30'b000000001000000000110011110000
                ;mem[1254] <= 30'b000000001000000000110100000000
                ;mem[1255] <= 30'b000000001000000000110100010000
                ;mem[1256] <= 30'b000000001000000000110111110000
                ;mem[1257] <= 30'b000000001000000000111000000000
                ;mem[1258] <= 30'b000000001000000000111000010000
                ;mem[1259] <= 30'b000000001000000000111000100000
                ;mem[1260] <= 30'b000000001000000000111000110000
                ;mem[1261] <= 30'b000000001000000000111001000000
                ;mem[1262] <= 30'b000000001000000000111001010000
                ;mem[1263] <= 30'b000000001000000000111001100000
                ;mem[1264] <= 30'b000000001000000000111001110000
                ;mem[1265] <= 30'b000000001000000000111010000000
                ;mem[1266] <= 30'b000000001000000000111010010000
                ;mem[1267] <= 30'b000000001000000000111010100000
                ;mem[1268] <= 30'b000000001000000000111010110000
                ;mem[1269] <= 30'b000000001000000000111011000000
                ;mem[1270] <= 30'b000000001000000000111111010000
                ;mem[1271] <= 30'b000000001000000000111111100000
                ;mem[1272] <= 30'b000000001000000000111111110000
                ;mem[1273] <= 30'b000000010000000000000000100000
                ;mem[1274] <= 30'b000000010000000000000000110000
                ;mem[1275] <= 30'b000000010000000000000001000000
                ;mem[1276] <= 30'b000000010000000000000001010000
                ;mem[1277] <= 30'b000000010000000000000001100000
                ;mem[1278] <= 30'b000000010000000000000100110000
                ;mem[1279] <= 30'b000000010000000000000101000000
                ;mem[1280] <= 30'b000000010000000000000101010000
                ;mem[1281] <= 30'b000000010000000000000101110000
                ;mem[1282] <= 30'b000000010000000000000110000000
                ;mem[1283] <= 30'b000000010000000000000110010000
                ;mem[1284] <= 30'b000000010000000000000110100000
                ;mem[1285] <= 30'b000000010000000000000110110000
                ;mem[1286] <= 30'b000000010000000000000111000000
                ;mem[1287] <= 30'b000000010000000000000111010000
                ;mem[1288] <= 30'b000000010000000000000111100000
                ;mem[1289] <= 30'b000000010000000000000111110000
                ;mem[1290] <= 30'b000000010000000000001000000000
                ;mem[1291] <= 30'b000000010000000000001000010000
                ;mem[1292] <= 30'b000000010000000000001011110000
                ;mem[1293] <= 30'b000000010000000000001100000000
                ;mem[1294] <= 30'b000000010000000000001100010000
                ;mem[1295] <= 30'b000000010000000000001100100000
                ;mem[1296] <= 30'b000000010000000000001100110000
                ;mem[1297] <= 30'b000000010000000000001101000000
                ;mem[1298] <= 30'b000000010000000000001101010000
                ;mem[1299] <= 30'b000000010000000000001101100000
                ;mem[1300] <= 30'b000000010000000000001101110000
                ;mem[1301] <= 30'b000000010000000000001110000000
                ;mem[1302] <= 30'b000000010000000000001110010000
                ;mem[1303] <= 30'b000000010000000000001110100000
                ;mem[1304] <= 30'b000000010000000000001110110000
                ;mem[1305] <= 30'b000000010000000000001111000000
                ;mem[1306] <= 30'b000000010000000000010011010000
                ;mem[1307] <= 30'b000000010000000000010011100000
                ;mem[1308] <= 30'b000000010000000000010011110000
                ;mem[1309] <= 30'b000000010000000000010100000000
                ;mem[1310] <= 30'b000000010000000000010100010000
                ;mem[1311] <= 30'b000000010000000000010100100000
                ;mem[1312] <= 30'b000000010000000000010100110000
                ;mem[1313] <= 30'b000000010000000000010101000000
                ;mem[1314] <= 30'b000000010000000000010101010000
                ;mem[1315] <= 30'b000000010000000000010101100000
                ;mem[1316] <= 30'b000000010000000000010101110000
                ;mem[1317] <= 30'b000000010000000000011011100000
                ;mem[1318] <= 30'b000000010000000000011011110000
                ;mem[1319] <= 30'b000000010000000000011100000000
                ;mem[1320] <= 30'b000000010000000000011100010000
                ;mem[1321] <= 30'b000000010000000000100010100000
                ;mem[1322] <= 30'b000000010000000000100010110000
                ;mem[1323] <= 30'b000000010000000000100011000000
                ;mem[1324] <= 30'b000000010000000000101001010000
                ;mem[1325] <= 30'b000000010000000000101001100000
                ;mem[1326] <= 30'b000000010000000000101001110000
                ;mem[1327] <= 30'b000000010000000000101010000000
                ;mem[1328] <= 30'b000000010000000000110000000000
                ;mem[1329] <= 30'b000000010000000000110000010000
                ;mem[1330] <= 30'b000000010000000000110000100000
                ;mem[1331] <= 30'b000000010000000000110000110000
                ;mem[1332] <= 30'b000000010000000000110110110000
                ;mem[1333] <= 30'b000000010000000000110111000000
                ;mem[1334] <= 30'b000000010000000000110111010000
                ;mem[1335] <= 30'b000000010000000000110111100000
                ;mem[1336] <= 30'b000000010000000000111101110000
                ;mem[1337] <= 30'b000000010000000000111110000000
                ;mem[1338] <= 30'b000000010000000000111110010000
                ;mem[1339] <= 30'b000000010000000000111110100000
                ;mem[1340] <= 30'b000000000000000001000100000000
                ;mem[1341] <= 30'b000000000000000001000100010000
                ;mem[1342] <= 30'b000000000000000001000100100000
                ;mem[1343] <= 30'b000000000000000001000100110000
                ;mem[1344] <= 30'b000000000000000001001010110000
                ;mem[1345] <= 30'b000000000000000001001011000000
                ;mem[1346] <= 30'b000000000000000001001011010000
                ;mem[1347] <= 30'b000000000000000001001011100000
                ;mem[1348] <= 30'b000000000000000001010001110000
                ;mem[1349] <= 30'b000000000000000001010010000000
                ;mem[1350] <= 30'b000000000000000001010010010000
                ;mem[1351] <= 30'b000000000000000001010010100000
                ;mem[1352] <= 30'b000000000000000001011000100000
                ;mem[1353] <= 30'b000000000000000001011000110000
                ;mem[1354] <= 30'b000000000000000001011001000000
                ;mem[1355] <= 30'b000000000000000001011001010000
                ;mem[1356] <= 30'b000000000000000001011111100000
                ;mem[1357] <= 30'b000000000000000001011111110000
                ;mem[1358] <= 30'b000000000000000001100000000000
                ;mem[1359] <= 30'b000000000000000001100110010000
                ;mem[1360] <= 30'b000000000000000001100110100000
                ;mem[1361] <= 30'b000000000000000001100110110000
                ;mem[1362] <= 30'b000000000000000001100111000000
                ;mem[1363] <= 30'b000000000000000001101101010000
                ;mem[1364] <= 30'b000000000000000001101101100000
                ;mem[1365] <= 30'b000000000000000001101101110000
                ;mem[1366] <= 30'b000000000000000001110100100000
                ;mem[1367] <= 30'b000000000000000000011111110000
                ;mem[1368] <= 30'b000000000000000000100101100000
                ;mem[1369] <= 30'b000000000000000000100101110000
                ;mem[1370] <= 30'b000000000000000000100110000000
                ;mem[1371] <= 30'b000000000000000000100110010000
                ;mem[1372] <= 30'b000000000000000000100110100000
                ;mem[1373] <= 30'b000000000000000000100110110000
                ;mem[1374] <= 30'b000000000000000000100111000000
                ;mem[1375] <= 30'b000000000000000000100111010000
                ;mem[1376] <= 30'b000000000000000000100111100000
                ;mem[1377] <= 30'b000000000000000000100111110000
                ;mem[1378] <= 30'b000000000000000000101100010000
                ;mem[1379] <= 30'b000000000000000000101100100000
                ;mem[1380] <= 30'b000000000000000000101100110000
                ;mem[1381] <= 30'b000000000000000000101101000000
                ;mem[1382] <= 30'b000000000000000000101101010000
                ;mem[1383] <= 30'b000000000000000000101101100000
                ;mem[1384] <= 30'b000000000000000000101101110000
                ;mem[1385] <= 30'b000000000000000000101110000000
                ;mem[1386] <= 30'b000000000000000000101110010000
                ;mem[1387] <= 30'b000000000000000000101110100000
                ;mem[1388] <= 30'b000000000000000000101110110000
                ;mem[1389] <= 30'b000000000000000000101111000000
                ;mem[1390] <= 30'b000000000000000000110011010000
                ;mem[1391] <= 30'b000000000000000000110011100000
                ;mem[1392] <= 30'b000000000000000000110011110000
                ;mem[1393] <= 30'b000000000000000000110101100000
                ;mem[1394] <= 30'b000000000000000000110101110000
                ;mem[1395] <= 30'b000000000000000000110110000000
                ;mem[1396] <= 30'b000000000000000000110110010000
                ;mem[1397] <= 30'b000000000000000000111010010000
                ;mem[1398] <= 30'b000000000000000000111010100000
                ;mem[1399] <= 30'b000000000000000000111100110000
                ;mem[1400] <= 30'b000000000000000000111101000000
                ;mem[1401] <= 30'b000000000000000000111101010000
                ;mem[1402] <= 30'b000000001000000000000000010000
                ;mem[1403] <= 30'b000000001000000000000000100000
                ;mem[1404] <= 30'b000000001000000000000000110000
                ;mem[1405] <= 30'b000000001000000000000001000000
                ;mem[1406] <= 30'b000000001000000000000001010000
                ;mem[1407] <= 30'b000000001000000000000001100000
                ;mem[1408] <= 30'b000000001000000000000001110000
                ;mem[1409] <= 30'b000000001000000000000010000000
                ;mem[1410] <= 30'b000000001000000000000010010000
                ;mem[1411] <= 30'b000000001000000000000010100000
                ;mem[1412] <= 30'b000000001000000000000010110000
                ;mem[1413] <= 30'b000000001000000000000011000000
                ;mem[1414] <= 30'b000000001000000000000111010000
                ;mem[1415] <= 30'b000000001000000000000111100000
                ;mem[1416] <= 30'b000000001000000000000111110000
                ;mem[1417] <= 30'b000000001000000000001001100000
                ;mem[1418] <= 30'b000000001000000000001001110000
                ;mem[1419] <= 30'b000000001000000000001010000000
                ;mem[1420] <= 30'b000000001000000000001010010000
                ;mem[1421] <= 30'b000000001000000000001110010000
                ;mem[1422] <= 30'b000000001000000000001110100000
                ;mem[1423] <= 30'b000000001000000000010000110000
                ;mem[1424] <= 30'b000000001000000000010001000000
                ;mem[1425] <= 30'b000000001000000000010001010000
                ;mem[1426] <= 30'b000000001000000000010101010000
                ;mem[1427] <= 30'b000000001000000000010101100000
                ;mem[1428] <= 30'b000000001000000000011000000000
                ;mem[1429] <= 30'b000000001000000000011000010000
                ;mem[1430] <= 30'b000000001000000000011000100000
                ;mem[1431] <= 30'b000000001000000000011100000000
                ;mem[1432] <= 30'b000000001000000000011100010000
                ;mem[1433] <= 30'b000000001000000000011111000000
                ;mem[1434] <= 30'b000000001000000000011111010000
                ;mem[1435] <= 30'b000000001000000000011111100000
                ;mem[1436] <= 30'b000000001000000000100011000000
                ;mem[1437] <= 30'b000000001000000000100011010000
                ;mem[1438] <= 30'b000000001000000000100110010000
                ;mem[1439] <= 30'b000000001000000000100110100000
                ;mem[1440] <= 30'b000000001000000000101010000000
                ;mem[1441] <= 30'b000000001000000000101010010000
                ;mem[1442] <= 30'b000000001000000000101101010000
                ;mem[1443] <= 30'b000000001000000000101101100000
                ;mem[1444] <= 30'b000000001000000000110000110000
                ;mem[1445] <= 30'b000000001000000000110001000000
                ;mem[1446] <= 30'b000000001000000000110100010000
                ;mem[1447] <= 30'b000000001000000000110100100000
                ;mem[1448] <= 30'b000000001000000000110111110000
                ;mem[1449] <= 30'b000000001000000000111000000000
                ;mem[1450] <= 30'b000000001000000000111011010000
                ;mem[1451] <= 30'b000000001000000000111011100000
                ;mem[1452] <= 30'b000000001000000000111110110000
                ;mem[1453] <= 30'b000000001000000000111111000000
                ;mem[1454] <= 30'b000000010000000000000001010000
                ;mem[1455] <= 30'b000000010000000000000001100000
                ;mem[1456] <= 30'b000000010000000000000100110000
                ;mem[1457] <= 30'b000000010000000000000101000000
                ;mem[1458] <= 30'b000000010000000000001000010000
                ;mem[1459] <= 30'b000000010000000000001000100000
                ;mem[1460] <= 30'b000000010000000000001011110000
                ;mem[1461] <= 30'b000000010000000000001100000000
                ;mem[1462] <= 30'b000000010000000000001111010000
                ;mem[1463] <= 30'b000000010000000000001111100000
                ;mem[1464] <= 30'b000000010000000000010010110000
                ;mem[1465] <= 30'b000000010000000000010011000000
                ;mem[1466] <= 30'b000000010000000000010110010000
                ;mem[1467] <= 30'b000000010000000000010110100000
                ;mem[1468] <= 30'b000000010000000000011001110000
                ;mem[1469] <= 30'b000000010000000000011010000000
                ;mem[1470] <= 30'b000000010000000000011101000000
                ;mem[1471] <= 30'b000000010000000000011101010000
                ;mem[1472] <= 30'b000000010000000000011101100000
                ;mem[1473] <= 30'b000000010000000000100000110000
                ;mem[1474] <= 30'b000000010000000000100001000000
                ;mem[1475] <= 30'b000000010000000000100100000000
                ;mem[1476] <= 30'b000000010000000000100100010000
                ;mem[1477] <= 30'b000000010000000000100111110000
                ;mem[1478] <= 30'b000000010000000000101000000000
                ;mem[1479] <= 30'b000000010000000000101010110000
                ;mem[1480] <= 30'b000000010000000000101011000000
                ;mem[1481] <= 30'b000000010000000000101011010000
                ;mem[1482] <= 30'b000000010000000000101110110000
                ;mem[1483] <= 30'b000000010000000000101111000000
                ;mem[1484] <= 30'b000000010000000000110001100000
                ;mem[1485] <= 30'b000000010000000000110001110000
                ;mem[1486] <= 30'b000000010000000000110010000000
                ;mem[1487] <= 30'b000000010000000000110101110000
                ;mem[1488] <= 30'b000000010000000000110110000000
                ;mem[1489] <= 30'b000000010000000000111000000000
                ;mem[1490] <= 30'b000000010000000000111000010000
                ;mem[1491] <= 30'b000000010000000000111000100000
                ;mem[1492] <= 30'b000000010000000000111000110000
                ;mem[1493] <= 30'b000000010000000000111100110000
                ;mem[1494] <= 30'b000000010000000000111101000000
                ;mem[1495] <= 30'b000000010000000000111101010000
                ;mem[1496] <= 30'b000000010000000000111101100000
                ;mem[1497] <= 30'b000000010000000000111101110000
                ;mem[1498] <= 30'b000000010000000000111110000000
                ;mem[1499] <= 30'b000000010000000000111110010000
                ;mem[1500] <= 30'b000000010000000000111110100000
                ;mem[1501] <= 30'b000000010000000000111110110000
                ;mem[1502] <= 30'b000000010000000000111111000000
                ;mem[1503] <= 30'b000000010000000000111111010000
                ;mem[1504] <= 30'b000000010000000000111111100000
                ;mem[1505] <= 30'b000000010000000000111111110000
                ;mem[1506] <= 30'b000000000000000001000010110000
                ;mem[1507] <= 30'b000000000000000001000011000000
                ;mem[1508] <= 30'b000000000000000001000101100000
                ;mem[1509] <= 30'b000000000000000001000101110000
                ;mem[1510] <= 30'b000000000000000001000110000000
                ;mem[1511] <= 30'b000000000000000001001001110000
                ;mem[1512] <= 30'b000000000000000001001010000000
                ;mem[1513] <= 30'b000000000000000001001100000000
                ;mem[1514] <= 30'b000000000000000001001100010000
                ;mem[1515] <= 30'b000000000000000001001100100000
                ;mem[1516] <= 30'b000000000000000001001100110000
                ;mem[1517] <= 30'b000000000000000001010000110000
                ;mem[1518] <= 30'b000000000000000001010001000000
                ;mem[1519] <= 30'b000000000000000001010001010000
                ;mem[1520] <= 30'b000000000000000001010001100000
                ;mem[1521] <= 30'b000000000000000001010001110000
                ;mem[1522] <= 30'b000000000000000001010010000000
                ;mem[1523] <= 30'b000000000000000001010010010000
                ;mem[1524] <= 30'b000000000000000001010010100000
                ;mem[1525] <= 30'b000000000000000001010010110000
                ;mem[1526] <= 30'b000000000000000001010011000000
                ;mem[1527] <= 30'b000000000000000001010011010000
                ;mem[1528] <= 30'b000000000000000001010011100000
                ;mem[1529] <= 30'b000000000000000001010011110000
                ;mem[1530] <= 30'b000000000000000001011000000000
                ;mem[1531] <= 30'b000000000000000001011000010000
                ;mem[1532] <= 30'b000000000000000001011000100000
                ;mem[1533] <= 30'b000000000000000001011000110000
                ;mem[1534] <= 30'b000000000000000001011001000000
                ;mem[1535] <= 30'b000000000000000001011001010000
                ;mem[1536] <= 30'b000000000000000001011001100000
                ;mem[1537] <= 30'b000000000000000001011001110000
                ;mem[1538] <= 30'b000000000000000001011010000000
                ;mem[1539] <= 30'b000000000000000001011010010000
                ;mem[1540] <= 30'b000000000000000001011111010000
                ;mem[1541] <= 30'b000000000000000001011111100000
                ;mem[1542] <= 30'b000000000000000001011111110000
                ;mem[1543] <= 30'b000000000000000001100000000000
                ;mem[1544] <= 30'b000000000000000001100000010000
                ;mem[1545] <= 30'b000000000000000001100000100000
                ;mem[1546] <= 30'b000000000000000001100000110000
                ;mem[1547] <= 30'b000000000000000000010111110000
                ;mem[1548] <= 30'b000000000000000000011000000000
                ;mem[1549] <= 30'b000000000000000000011000010000
                ;mem[1550] <= 30'b000000000000000000011110100000
                ;mem[1551] <= 30'b000000000000000000011110110000
                ;mem[1552] <= 30'b000000000000000000011111000000
                ;mem[1553] <= 30'b000000000000000000100101100000
                ;mem[1554] <= 30'b000000000000000000100101110000
                ;mem[1555] <= 30'b000000000000000000101100010000
                ;mem[1556] <= 30'b000000000000000000101100100000
                ;mem[1557] <= 30'b000000000000000000110011010000
                ;mem[1558] <= 30'b000000000000000000110011100000
                ;mem[1559] <= 30'b000000000000000000111010010000
                ;mem[1560] <= 30'b000000000000000000111010100000
                ;mem[1561] <= 30'b000000001000000000000000010000
                ;mem[1562] <= 30'b000000001000000000000000100000
                ;mem[1563] <= 30'b000000001000000000000111010000
                ;mem[1564] <= 30'b000000001000000000000111100000
                ;mem[1565] <= 30'b000000001000000000001110010000
                ;mem[1566] <= 30'b000000001000000000001110100000
                ;mem[1567] <= 30'b000000001000000000010101000000
                ;mem[1568] <= 30'b000000001000000000010101010000
                ;mem[1569] <= 30'b000000001000000000010101100000
                ;mem[1570] <= 30'b000000001000000000011100000000
                ;mem[1571] <= 30'b000000001000000000011100010000
                ;mem[1572] <= 30'b000000001000000000011110000000
                ;mem[1573] <= 30'b000000001000000000011110010000
                ;mem[1574] <= 30'b000000001000000000011110100000
                ;mem[1575] <= 30'b000000001000000000011110110000
                ;mem[1576] <= 30'b000000001000000000011111000000
                ;mem[1577] <= 30'b000000001000000000011111010000
                ;mem[1578] <= 30'b000000001000000000100011000000
                ;mem[1579] <= 30'b000000001000000000100011010000
                ;mem[1580] <= 30'b000000001000000000100100110000
                ;mem[1581] <= 30'b000000001000000000100101000000
                ;mem[1582] <= 30'b000000001000000000100101010000
                ;mem[1583] <= 30'b000000001000000000100101100000
                ;mem[1584] <= 30'b000000001000000000100101110000
                ;mem[1585] <= 30'b000000001000000000100110000000
                ;mem[1586] <= 30'b000000001000000000100110010000
                ;mem[1587] <= 30'b000000001000000000100110100000
                ;mem[1588] <= 30'b000000001000000000101010000000
                ;mem[1589] <= 30'b000000001000000000101010010000
                ;mem[1590] <= 30'b000000001000000000101011010000
                ;mem[1591] <= 30'b000000001000000000101011100000
                ;mem[1592] <= 30'b000000001000000000101011110000
                ;mem[1593] <= 30'b000000001000000000101100000000
                ;mem[1594] <= 30'b000000001000000000101100010000
                ;mem[1595] <= 30'b000000001000000000101101010000
                ;mem[1596] <= 30'b000000001000000000101101100000
                ;mem[1597] <= 30'b000000001000000000110000110000
                ;mem[1598] <= 30'b000000001000000000110001000000
                ;mem[1599] <= 30'b000000001000000000110010000000
                ;mem[1600] <= 30'b000000001000000000110010010000
                ;mem[1601] <= 30'b000000001000000000110010100000
                ;mem[1602] <= 30'b000000001000000000110010110000
                ;mem[1603] <= 30'b000000001000000000110100010000
                ;mem[1604] <= 30'b000000001000000000110100100000
                ;mem[1605] <= 30'b000000001000000000110111110000
                ;mem[1606] <= 30'b000000001000000000111000000000
                ;mem[1607] <= 30'b000000001000000000111001000000
                ;mem[1608] <= 30'b000000001000000000111001010000
                ;mem[1609] <= 30'b000000001000000000111001100000
                ;mem[1610] <= 30'b000000001000000000111011010000
                ;mem[1611] <= 30'b000000001000000000111011100000
                ;mem[1612] <= 30'b000000001000000000111110110000
                ;mem[1613] <= 30'b000000001000000000111111000000
                ;mem[1614] <= 30'b000000001000000000111111110000
                ;mem[1615] <= 30'b000000010000000000000000000000
                ;mem[1616] <= 30'b000000010000000000000000010000
                ;mem[1617] <= 30'b000000010000000000000001010000
                ;mem[1618] <= 30'b000000010000000000000001100000
                ;mem[1619] <= 30'b000000010000000000000100110000
                ;mem[1620] <= 30'b000000010000000000000101000000
                ;mem[1621] <= 30'b000000010000000000000110000000
                ;mem[1622] <= 30'b000000010000000000000110010000
                ;mem[1623] <= 30'b000000010000000000000110100000
                ;mem[1624] <= 30'b000000010000000000000110110000
                ;mem[1625] <= 30'b000000010000000000001000010000
                ;mem[1626] <= 30'b000000010000000000001000100000
                ;mem[1627] <= 30'b000000010000000000001011110000
                ;mem[1628] <= 30'b000000010000000000001100000000
                ;mem[1629] <= 30'b000000010000000000001101000000
                ;mem[1630] <= 30'b000000010000000000001101010000
                ;mem[1631] <= 30'b000000010000000000001101100000
                ;mem[1632] <= 30'b000000010000000000001111010000
                ;mem[1633] <= 30'b000000010000000000001111100000
                ;mem[1634] <= 30'b000000010000000000010010110000
                ;mem[1635] <= 30'b000000010000000000010011000000
                ;mem[1636] <= 30'b000000010000000000010011110000
                ;mem[1637] <= 30'b000000010000000000010100000000
                ;mem[1638] <= 30'b000000010000000000010100010000
                ;mem[1639] <= 30'b000000010000000000010110010000
                ;mem[1640] <= 30'b000000010000000000010110100000
                ;mem[1641] <= 30'b000000010000000000011001110000
                ;mem[1642] <= 30'b000000010000000000011010000000
                ;mem[1643] <= 30'b000000010000000000011010110000
                ;mem[1644] <= 30'b000000010000000000011011000000
                ;mem[1645] <= 30'b000000010000000000011011010000
                ;mem[1646] <= 30'b000000010000000000011101010000
                ;mem[1647] <= 30'b000000010000000000011101100000
                ;mem[1648] <= 30'b000000010000000000100000110000
                ;mem[1649] <= 30'b000000010000000000100001000000
                ;mem[1650] <= 30'b000000010000000000100010000000
                ;mem[1651] <= 30'b000000010000000000100010010000
                ;mem[1652] <= 30'b000000010000000000100100000000
                ;mem[1653] <= 30'b000000010000000000100100010000
                ;mem[1654] <= 30'b000000010000000000100111110000
                ;mem[1655] <= 30'b000000010000000000101000000000
                ;mem[1656] <= 30'b000000010000000000101001010000
                ;mem[1657] <= 30'b000000010000000000101001100000
                ;mem[1658] <= 30'b000000010000000000101001110000
                ;mem[1659] <= 30'b000000010000000000101010110000
                ;mem[1660] <= 30'b000000010000000000101011000000
                ;mem[1661] <= 30'b000000010000000000101110110000
                ;mem[1662] <= 30'b000000010000000000101111000000
                ;mem[1663] <= 30'b000000010000000000101111010000
                ;mem[1664] <= 30'b000000010000000000110001010000
                ;mem[1665] <= 30'b000000010000000000110001100000
                ;mem[1666] <= 30'b000000010000000000110001110000
                ;mem[1667] <= 30'b000000010000000000110110000000
                ;mem[1668] <= 30'b000000010000000000110110010000
                ;mem[1669] <= 30'b000000010000000000110110100000
                ;mem[1670] <= 30'b000000010000000000110111100000
                ;mem[1671] <= 30'b000000010000000000110111110000
                ;mem[1672] <= 30'b000000010000000000111000000000
                ;mem[1673] <= 30'b000000010000000000111000010000
                ;mem[1674] <= 30'b000000010000000000111000100000
                ;mem[1675] <= 30'b000000010000000000111101010000
                ;mem[1676] <= 30'b000000010000000000111101100000
                ;mem[1677] <= 30'b000000010000000000111101110000
                ;mem[1678] <= 30'b000000010000000000111110000000
                ;mem[1679] <= 30'b000000010000000000111110010000
                ;mem[1680] <= 30'b000000010000000000111110100000
                ;mem[1681] <= 30'b000000010000000000111110110000
                ;mem[1682] <= 30'b000000010000000000111111000000
                ;mem[1683] <= 30'b000000010000000000111111010000
                ;mem[1684] <= 30'b000000000000000001000010110000
                ;mem[1685] <= 30'b000000000000000001000011000000
                ;mem[1686] <= 30'b000000000000000001000011010000
                ;mem[1687] <= 30'b000000000000000001000101010000
                ;mem[1688] <= 30'b000000000000000001000101100000
                ;mem[1689] <= 30'b000000000000000001000101110000
                ;mem[1690] <= 30'b000000000000000001001010000000
                ;mem[1691] <= 30'b000000000000000001001010010000
                ;mem[1692] <= 30'b000000000000000001001010100000
                ;mem[1693] <= 30'b000000000000000001001011100000
                ;mem[1694] <= 30'b000000000000000001001011110000
                ;mem[1695] <= 30'b000000000000000001001100000000
                ;mem[1696] <= 30'b000000000000000001001100010000
                ;mem[1697] <= 30'b000000000000000001001100100000
                ;mem[1698] <= 30'b000000000000000001010001010000
                ;mem[1699] <= 30'b000000000000000001010001100000
                ;mem[1700] <= 30'b000000000000000001010001110000
                ;mem[1701] <= 30'b000000000000000001010010000000
                ;mem[1702] <= 30'b000000000000000001010010010000
                ;mem[1703] <= 30'b000000000000000001010010100000
                ;mem[1704] <= 30'b000000000000000001010010110000
                ;mem[1705] <= 30'b000000000000000001010011000000
                ;mem[1706] <= 30'b000000000000000001010011010000
                ;mem[1707] <= 30'b000000000000000001011000110000
                ;mem[1708] <= 30'b000000000000000001011001000000
                ;mem[1709] <= 30'b000000000000000001011001010000
                ;mem[1710] <= 30'b000000000000000001011001100000
                ;mem[1711] <= 30'b000000000000000001011001110000
                ;mem[1712] <= 30'b000000000000000000110100010000
                ;mem[1713] <= 30'b000000000000000000110100100000
                ;mem[1714] <= 30'b000000000000000000110100110000
                ;mem[1715] <= 30'b000000000000000000110101000000
                ;mem[1716] <= 30'b000000000000000000110101010000
                ;mem[1717] <= 30'b000000000000000000111011000000
                ;mem[1718] <= 30'b000000000000000000111011010000
                ;mem[1719] <= 30'b000000000000000000111011100000
                ;mem[1720] <= 30'b000000000000000000111011110000
                ;mem[1721] <= 30'b000000000000000000111100000000
                ;mem[1722] <= 30'b000000000000000000111100010000
                ;mem[1723] <= 30'b000000000000000000111100100000
                ;mem[1724] <= 30'b000000000000000000111100110000
                ;mem[1725] <= 30'b000000000000000000111101000000
                ;mem[1726] <= 30'b000000001000000000001000010000
                ;mem[1727] <= 30'b000000001000000000001000100000
                ;mem[1728] <= 30'b000000001000000000001000110000
                ;mem[1729] <= 30'b000000001000000000001001000000
                ;mem[1730] <= 30'b000000001000000000001001010000
                ;mem[1731] <= 30'b000000001000000000001111000000
                ;mem[1732] <= 30'b000000001000000000001111010000
                ;mem[1733] <= 30'b000000001000000000001111100000
                ;mem[1734] <= 30'b000000001000000000001111110000
                ;mem[1735] <= 30'b000000001000000000010000000000
                ;mem[1736] <= 30'b000000001000000000010000010000
                ;mem[1737] <= 30'b000000001000000000010000100000
                ;mem[1738] <= 30'b000000001000000000010000110000
                ;mem[1739] <= 30'b000000001000000000010001000000
                ;mem[1740] <= 30'b000000001000000000010101110000
                ;mem[1741] <= 30'b000000001000000000010110000000
                ;mem[1742] <= 30'b000000001000000000010110010000
                ;mem[1743] <= 30'b000000001000000000010111110000
                ;mem[1744] <= 30'b000000001000000000011000000000
                ;mem[1745] <= 30'b000000001000000000011100100000
                ;mem[1746] <= 30'b000000001000000000011100110000
                ;mem[1747] <= 30'b000000001000000000011101000000
                ;mem[1748] <= 30'b000000001000000000011110100000
                ;mem[1749] <= 30'b000000001000000000011110110000
                ;mem[1750] <= 30'b000000001000000000011111000000
                ;mem[1751] <= 30'b000000001000000000100011010000
                ;mem[1752] <= 30'b000000001000000000100011100000
                ;mem[1753] <= 30'b000000001000000000100011110000
                ;mem[1754] <= 30'b000000001000000000100101100000
                ;mem[1755] <= 30'b000000001000000000100101110000
                ;mem[1756] <= 30'b000000001000000000101010000000
                ;mem[1757] <= 30'b000000001000000000101010010000
                ;mem[1758] <= 30'b000000001000000000101010100000
                ;mem[1759] <= 30'b000000001000000000101100010000
                ;mem[1760] <= 30'b000000001000000000101100100000
                ;mem[1761] <= 30'b000000001000000000101100110000
                ;mem[1762] <= 30'b000000001000000000110001000000
                ;mem[1763] <= 30'b000000001000000000110001010000
                ;mem[1764] <= 30'b000000001000000000110001100000
                ;mem[1765] <= 30'b000000001000000000110011000000
                ;mem[1766] <= 30'b000000001000000000110011010000
                ;mem[1767] <= 30'b000000001000000000110011100000
                ;mem[1768] <= 30'b000000001000000000111000000000
                ;mem[1769] <= 30'b000000001000000000111000010000
                ;mem[1770] <= 30'b000000001000000000111000100000
                ;mem[1771] <= 30'b000000001000000000111001110000
                ;mem[1772] <= 30'b000000001000000000111010000000
                ;mem[1773] <= 30'b000000001000000000111010010000
                ;mem[1774] <= 30'b000000001000000000111010100000
                ;mem[1775] <= 30'b000000001000000000111111000000
                ;mem[1776] <= 30'b000000001000000000111111010000
                ;mem[1777] <= 30'b000000001000000000111111100000
                ;mem[1778] <= 30'b000000001000000000111111110000
                ;mem[1779] <= 30'b000000010000000000000000010000
                ;mem[1780] <= 30'b000000010000000000000000100000
                ;mem[1781] <= 30'b000000010000000000000000110000
                ;mem[1782] <= 30'b000000010000000000000101000000
                ;mem[1783] <= 30'b000000010000000000000101010000
                ;mem[1784] <= 30'b000000010000000000000101100000
                ;mem[1785] <= 30'b000000010000000000000111000000
                ;mem[1786] <= 30'b000000010000000000000111010000
                ;mem[1787] <= 30'b000000010000000000000111100000
                ;mem[1788] <= 30'b000000010000000000001100000000
                ;mem[1789] <= 30'b000000010000000000001100010000
                ;mem[1790] <= 30'b000000010000000000001100100000
                ;mem[1791] <= 30'b000000010000000000001101110000
                ;mem[1792] <= 30'b000000010000000000001110000000
                ;mem[1793] <= 30'b000000010000000000001110010000
                ;mem[1794] <= 30'b000000010000000000001110100000
                ;mem[1795] <= 30'b000000010000000000010011000000
                ;mem[1796] <= 30'b000000010000000000010011010000
                ;mem[1797] <= 30'b000000010000000000010011100000
                ;mem[1798] <= 30'b000000010000000000010011110000
                ;mem[1799] <= 30'b000000010000000000010100000000
                ;mem[1800] <= 30'b000000010000000000010100010000
                ;mem[1801] <= 30'b000000010000000000010100100000
                ;mem[1802] <= 30'b000000010000000000010100110000
                ;mem[1803] <= 30'b000000010000000000010101000000
                ;mem[1804] <= 30'b000000010000000000010101010000
                ;mem[1805] <= 30'b000000010000000000010101100000
                ;mem[1806] <= 30'b000000010000000000011010010000
                ;mem[1807] <= 30'b000000010000000000011010100000
                ;mem[1808] <= 30'b000000010000000000011010110000
                ;mem[1809] <= 30'b000000010000000000011011000000
                ;mem[1810] <= 30'b000000010000000000011011010000
                ;mem[1811] <= 30'b000000010000000000011011100000
                ;mem[1812] <= 30'b000000010000000000011100000000
                ;mem[1813] <= 30'b000000010000000000011100010000
                ;mem[1814] <= 30'b000000010000000000100010110000
                ;mem[1815] <= 30'b000000010000000000100011000000
                ;mem[1816] <= 30'b000000010000000000100011010000
                ;mem[1817] <= 30'b000000010000000000101001110000
                ;mem[1818] <= 30'b000000010000000000101010000000
                ;mem[1819] <= 30'b000000010000000000101010010000
                ;mem[1820] <= 30'b000000010000000000110000110000
                ;mem[1821] <= 30'b000000010000000000110001000000
                ;mem[1822] <= 30'b000000010000000000110111100000
                ;mem[1823] <= 30'b000000010000000000110111110000
                ;mem[1824] <= 30'b000000010000000000111000000000
                ;mem[1825] <= 30'b000000010000000000111110100000
                ;mem[1826] <= 30'b000000010000000000111110110000
                ;mem[1827] <= 30'b000000000000000001000100110000
                ;mem[1828] <= 30'b000000000000000001000101000000
                ;mem[1829] <= 30'b000000000000000001001011100000
                ;mem[1830] <= 30'b000000000000000001001011110000
                ;mem[1831] <= 30'b000000000000000001001100000000
                ;mem[1832] <= 30'b000000000000000001010010100000
                ;mem[1833] <= 30'b000000000000000001010010110000
                ;mem[1834] <= 30'b000000000000000001011001100000
                ;mem[1835] <= 30'b000000000000000001011001110000
                ;mem[1836] <= 30'b000000000000000001100000100000
                ;mem[1837] <= 30'b000000000000000001100000110000
                ;mem[1838] <= 30'b000000000000000001100111010000
                ;mem[1839] <= 30'b000000000000000001100111100000
                ;mem[1840] <= 30'b000000000000000001101110010000
                ;mem[1841] <= 30'b000000000000000001101110100000
                ;mem[1842] <= 30'b000000000000000001110101100000
                ;mem[1843] <= 30'b000000000000000000100110100000
                ;mem[1844] <= 30'b000000000000000000100110110000
                ;mem[1845] <= 30'b000000000000000000100111000000
                ;mem[1846] <= 30'b000000000000000000100111010000
                ;mem[1847] <= 30'b000000000000000000100111100000
                ;mem[1848] <= 30'b000000000000000000101101000000
                ;mem[1849] <= 30'b000000000000000000101101010000
                ;mem[1850] <= 30'b000000000000000000101101100000
                ;mem[1851] <= 30'b000000000000000000101101110000
                ;mem[1852] <= 30'b000000000000000000101110000000
                ;mem[1853] <= 30'b000000000000000000101110010000
                ;mem[1854] <= 30'b000000000000000000101110100000
                ;mem[1855] <= 30'b000000000000000000101110110000
                ;mem[1856] <= 30'b000000000000000000110011110000
                ;mem[1857] <= 30'b000000000000000000110100000000
                ;mem[1858] <= 30'b000000000000000000110100010000
                ;mem[1859] <= 30'b000000000000000000110100100000
                ;mem[1860] <= 30'b000000000000000000110100110000
                ;mem[1861] <= 30'b000000000000000000110101000000
                ;mem[1862] <= 30'b000000000000000000110101010000
                ;mem[1863] <= 30'b000000000000000000110101100000
                ;mem[1864] <= 30'b000000000000000000110101110000
                ;mem[1865] <= 30'b000000000000000000111010100000
                ;mem[1866] <= 30'b000000000000000000111010110000
                ;mem[1867] <= 30'b000000000000000000111011000000
                ;mem[1868] <= 30'b000000000000000000111011010000
                ;mem[1869] <= 30'b000000000000000000111100000000
                ;mem[1870] <= 30'b000000000000000000111100010000
                ;mem[1871] <= 30'b000000000000000000111100100000
                ;mem[1872] <= 30'b000000000000000000111100110000
                ;mem[1873] <= 30'b000000001000000000000001000000
                ;mem[1874] <= 30'b000000001000000000000001010000
                ;mem[1875] <= 30'b000000001000000000000001100000
                ;mem[1876] <= 30'b000000001000000000000001110000
                ;mem[1877] <= 30'b000000001000000000000010000000
                ;mem[1878] <= 30'b000000001000000000000010010000
                ;mem[1879] <= 30'b000000001000000000000010100000
                ;mem[1880] <= 30'b000000001000000000000010110000
                ;mem[1881] <= 30'b000000001000000000000111110000
                ;mem[1882] <= 30'b000000001000000000001000000000
                ;mem[1883] <= 30'b000000001000000000001000010000
                ;mem[1884] <= 30'b000000001000000000001000100000
                ;mem[1885] <= 30'b000000001000000000001000110000
                ;mem[1886] <= 30'b000000001000000000001001000000
                ;mem[1887] <= 30'b000000001000000000001001010000
                ;mem[1888] <= 30'b000000001000000000001001100000
                ;mem[1889] <= 30'b000000001000000000001001110000
                ;mem[1890] <= 30'b000000001000000000001110100000
                ;mem[1891] <= 30'b000000001000000000001110110000
                ;mem[1892] <= 30'b000000001000000000001111000000
                ;mem[1893] <= 30'b000000001000000000001111010000
                ;mem[1894] <= 30'b000000001000000000010000000000
                ;mem[1895] <= 30'b000000001000000000010000010000
                ;mem[1896] <= 30'b000000001000000000010000100000
                ;mem[1897] <= 30'b000000001000000000010000110000
                ;mem[1898] <= 30'b000000001000000000010101010000
                ;mem[1899] <= 30'b000000001000000000010101100000
                ;mem[1900] <= 30'b000000001000000000010101110000
                ;mem[1901] <= 30'b000000001000000000010110000000
                ;mem[1902] <= 30'b000000001000000000010111100000
                ;mem[1903] <= 30'b000000001000000000010111110000
                ;mem[1904] <= 30'b000000001000000000011000000000
                ;mem[1905] <= 30'b000000001000000000011100010000
                ;mem[1906] <= 30'b000000001000000000011100100000
                ;mem[1907] <= 30'b000000001000000000011100110000
                ;mem[1908] <= 30'b000000001000000000011110100000
                ;mem[1909] <= 30'b000000001000000000011110110000
                ;mem[1910] <= 30'b000000001000000000011111000000
                ;mem[1911] <= 30'b000000001000000000011111010000
                ;mem[1912] <= 30'b000000001000000000100011000000
                ;mem[1913] <= 30'b000000001000000000100011010000
                ;mem[1914] <= 30'b000000001000000000100011100000
                ;mem[1915] <= 30'b000000001000000000100011110000
                ;mem[1916] <= 30'b000000001000000000100101110000
                ;mem[1917] <= 30'b000000001000000000100110000000
                ;mem[1918] <= 30'b000000001000000000100110010000
                ;mem[1919] <= 30'b000000001000000000101010000000
                ;mem[1920] <= 30'b000000001000000000101010010000
                ;mem[1921] <= 30'b000000001000000000101010100000
                ;mem[1922] <= 30'b000000001000000000101101000000
                ;mem[1923] <= 30'b000000001000000000101101010000
                ;mem[1924] <= 30'b000000001000000000110001000000
                ;mem[1925] <= 30'b000000001000000000110001010000
                ;mem[1926] <= 30'b000000001000000000110001100000
                ;mem[1927] <= 30'b000000001000000000110100000000
                ;mem[1928] <= 30'b000000001000000000110100010000
                ;mem[1929] <= 30'b000000001000000000111000000000
                ;mem[1930] <= 30'b000000001000000000111000010000
                ;mem[1931] <= 30'b000000001000000000111011000000
                ;mem[1932] <= 30'b000000001000000000111011010000
                ;mem[1933] <= 30'b000000001000000000111110110000
                ;mem[1934] <= 30'b000000001000000000111111000000
                ;mem[1935] <= 30'b000000001000000000111111010000
                ;mem[1936] <= 30'b000000010000000000000001000000
                ;mem[1937] <= 30'b000000010000000000000001010000
                ;mem[1938] <= 30'b000000010000000000000101000000
                ;mem[1939] <= 30'b000000010000000000000101010000
                ;mem[1940] <= 30'b000000010000000000000101100000
                ;mem[1941] <= 30'b000000010000000000001000000000
                ;mem[1942] <= 30'b000000010000000000001000010000
                ;mem[1943] <= 30'b000000010000000000001100000000
                ;mem[1944] <= 30'b000000010000000000001100010000
                ;mem[1945] <= 30'b000000010000000000001111000000
                ;mem[1946] <= 30'b000000010000000000001111010000
                ;mem[1947] <= 30'b000000010000000000010010110000
                ;mem[1948] <= 30'b000000010000000000010011000000
                ;mem[1949] <= 30'b000000010000000000010011010000
                ;mem[1950] <= 30'b000000010000000000010110000000
                ;mem[1951] <= 30'b000000010000000000010110010000
                ;mem[1952] <= 30'b000000010000000000011001110000
                ;mem[1953] <= 30'b000000010000000000011010000000
                ;mem[1954] <= 30'b000000010000000000011010010000
                ;mem[1955] <= 30'b000000010000000000011101000000
                ;mem[1956] <= 30'b000000010000000000011101010000
                ;mem[1957] <= 30'b000000010000000000100000110000
                ;mem[1958] <= 30'b000000010000000000100001000000
                ;mem[1959] <= 30'b000000010000000000100001010000
                ;mem[1960] <= 30'b000000010000000000100100000000
                ;mem[1961] <= 30'b000000010000000000100100010000
                ;mem[1962] <= 30'b000000010000000000100111110000
                ;mem[1963] <= 30'b000000010000000000101000000000
                ;mem[1964] <= 30'b000000010000000000101000010000
                ;mem[1965] <= 30'b000000010000000000101010110000
                ;mem[1966] <= 30'b000000010000000000101011000000
                ;mem[1967] <= 30'b000000010000000000101111000000
                ;mem[1968] <= 30'b000000010000000000101111010000
                ;mem[1969] <= 30'b000000010000000000101111100000
                ;mem[1970] <= 30'b000000010000000000110001110000
                ;mem[1971] <= 30'b000000010000000000110010000000
                ;mem[1972] <= 30'b000000010000000000110110010000
                ;mem[1973] <= 30'b000000010000000000110110100000
                ;mem[1974] <= 30'b000000010000000000111000100000
                ;mem[1975] <= 30'b000000010000000000111000110000
                ;mem[1976] <= 30'b000000010000000000111001000000
                ;mem[1977] <= 30'b000000010000000000111101010000
                ;mem[1978] <= 30'b000000010000000000111101100000
                ;mem[1979] <= 30'b000000010000000000111111100000
                ;mem[1980] <= 30'b000000010000000000111111110000
                ;mem[1981] <= 30'b000000000000000001000011000000
                ;mem[1982] <= 30'b000000000000000001000011010000
                ;mem[1983] <= 30'b000000000000000001000011100000
                ;mem[1984] <= 30'b000000000000000001000101110000
                ;mem[1985] <= 30'b000000000000000001000110000000
                ;mem[1986] <= 30'b000000000000000001001010010000
                ;mem[1987] <= 30'b000000000000000001001010100000
                ;mem[1988] <= 30'b000000000000000001001100100000
                ;mem[1989] <= 30'b000000000000000001001100110000
                ;mem[1990] <= 30'b000000000000000001001101000000
                ;mem[1991] <= 30'b000000000000000001010001010000
                ;mem[1992] <= 30'b000000000000000001010001100000
                ;mem[1993] <= 30'b000000000000000001010011100000
                ;mem[1994] <= 30'b000000000000000001010011110000
                ;mem[1995] <= 30'b000000000000000001011000100000
                ;mem[1996] <= 30'b000000000000000001011000110000
                ;mem[1997] <= 30'b000000000000000001011001000000
                ;mem[1998] <= 30'b000000000000000001011010010000
                ;mem[1999] <= 30'b000000000000000001011010100000
                ;mem[2000] <= 30'b000000000000000001011010110000
                ;mem[2001] <= 30'b000000000000000001011111110000
                ;mem[2002] <= 30'b000000000000000001100000000000
                ;mem[2003] <= 30'b000000000000000001100000010000
                ;mem[2004] <= 30'b000000000000000001100000110000
                ;mem[2005] <= 30'b000000000000000001100001000000
                ;mem[2006] <= 30'b000000000000000001100001010000
                ;mem[2007] <= 30'b000000000000000001100001100000
                ;mem[2008] <= 30'b000000000000000001100111010000
                ;mem[2009] <= 30'b000000000000000001100111100000
                ;mem[2010] <= 30'b000000000000000001100111110000
                ;mem[2011] <= 30'b000000000000000001101000000000
                ;mem[2012] <= 30'b000000000000000000011111010000
                ;mem[2013] <= 30'b000000000000000000011111100000
                ;mem[2014] <= 30'b000000000000000000011111110000
                ;mem[2015] <= 30'b000000000000000000100110010000
                ;mem[2016] <= 30'b000000000000000000100110100000
                ;mem[2017] <= 30'b000000000000000000100110110000
                ;mem[2018] <= 30'b000000000000000000101101010000
                ;mem[2019] <= 30'b000000000000000000101101100000
                ;mem[2020] <= 30'b000000000000000000101101110000
                ;mem[2021] <= 30'b000000000000000000101110000000
                ;mem[2022] <= 30'b000000000000000000110100010000
                ;mem[2023] <= 30'b000000000000000000110100100000
                ;mem[2024] <= 30'b000000000000000000110100110000
                ;mem[2025] <= 30'b000000000000000000111011010000
                ;mem[2026] <= 30'b000000000000000000111011100000
                ;mem[2027] <= 30'b000000000000000000111011110000
                ;mem[2028] <= 30'b000000001000000000000001010000
                ;mem[2029] <= 30'b000000001000000000000001100000
                ;mem[2030] <= 30'b000000001000000000000001110000
                ;mem[2031] <= 30'b000000001000000000000010000000
                ;mem[2032] <= 30'b000000001000000000001000010000
                ;mem[2033] <= 30'b000000001000000000001000100000
                ;mem[2034] <= 30'b000000001000000000001000110000
                ;mem[2035] <= 30'b000000001000000000001111010000
                ;mem[2036] <= 30'b000000001000000000001111100000
                ;mem[2037] <= 30'b000000001000000000001111110000
                ;mem[2038] <= 30'b000000001000000000010110010000
                ;mem[2039] <= 30'b000000001000000000010110100000
                ;mem[2040] <= 30'b000000001000000000010110110000
                ;mem[2041] <= 30'b000000001000000000010111000000
                ;mem[2042] <= 30'b000000001000000000011101010000
                ;mem[2043] <= 30'b000000001000000000011101100000
                ;mem[2044] <= 30'b000000001000000000011101110000
                ;mem[2045] <= 30'b000000001000000000011110000000
                ;mem[2046] <= 30'b000000001000000000100100010000
                ;mem[2047] <= 30'b000000001000000000100100100000
                ;mem[2048] <= 30'b000000001000000000100100110000
                ;mem[2049] <= 30'b000000001000000000100101000000
                ;mem[2050] <= 30'b000000001000000000101011010000
                ;mem[2051] <= 30'b000000001000000000101011100000
                ;mem[2052] <= 30'b000000001000000000101011110000
                ;mem[2053] <= 30'b000000001000000000101100000000
                ;mem[2054] <= 30'b000000001000000000110010010000
                ;mem[2055] <= 30'b000000001000000000110010100000
                ;mem[2056] <= 30'b000000001000000000110010110000
                ;mem[2057] <= 30'b000000001000000000110011000000
                ;mem[2058] <= 30'b000000001000000000111001010000
                ;mem[2059] <= 30'b000000001000000000111001100000
                ;mem[2060] <= 30'b000000001000000000111001110000
                ;mem[2061] <= 30'b000000010000000000000000000000
                ;mem[2062] <= 30'b000000010000000000000110010000
                ;mem[2063] <= 30'b000000010000000000000110100000
                ;mem[2064] <= 30'b000000010000000000000110110000
                ;mem[2065] <= 30'b000000010000000000000111000000
                ;mem[2066] <= 30'b000000010000000000001101010000
                ;mem[2067] <= 30'b000000010000000000001101100000
                ;mem[2068] <= 30'b000000010000000000001101110000
                ;mem[2069] <= 30'b000000010000000000010100010000
                ;mem[2070] <= 30'b000000010000000000010100100000
                ;mem[2071] <= 30'b000000010000000000010100110000
                ;mem[2072] <= 30'b000000010000000000011011010000
                ;mem[2073] <= 30'b000000010000000000011011100000
                ;mem[2074] <= 30'b000000010000000000011011110000
                ;mem[2075] <= 30'b000000010000000000100010010000
                ;mem[2076] <= 30'b000000010000000000100010100000
                ;mem[2077] <= 30'b000000010000000000100010110000
                ;mem[2078] <= 30'b000000010000000000101001010000
                ;mem[2079] <= 30'b000000010000000000101001100000
                ;mem[2080] <= 30'b000000010000000000101001110000
                ;mem[2081] <= 30'b000000010000000000101010000000
                ;mem[2082] <= 30'b000000010000000000110000010000
                ;mem[2083] <= 30'b000000010000000000110000100000
                ;mem[2084] <= 30'b000000010000000000110000110000
                ;mem[2085] <= 30'b000000010000000000110001000000
                ;mem[2086] <= 30'b000000010000000000110111010000
                ;mem[2087] <= 30'b000000010000000000110111100000
                ;mem[2088] <= 30'b000000010000000000110111110000
                ;mem[2089] <= 30'b000000010000000000111000000000
                ;mem[2090] <= 30'b000000010000000000111110000000
                ;mem[2091] <= 30'b000000010000000000111110010000
                ;mem[2092] <= 30'b000000010000000000111110100000
                ;mem[2093] <= 30'b000000010000000000111110110000
                ;mem[2094] <= 30'b000000010000000000111111000000
                ;mem[2095] <= 30'b000000000000000001000100010000
                ;mem[2096] <= 30'b000000000000000001000100100000
                ;mem[2097] <= 30'b000000000000000001000100110000
                ;mem[2098] <= 30'b000000000000000001000101000000
                ;mem[2099] <= 30'b000000000000000001001011010000
                ;mem[2100] <= 30'b000000000000000001001011100000
                ;mem[2101] <= 30'b000000000000000001001011110000
                ;mem[2102] <= 30'b000000000000000001001100000000
                ;mem[2103] <= 30'b000000000000000001010010000000
                ;mem[2104] <= 30'b000000000000000001010010010000
                ;mem[2105] <= 30'b000000000000000001010010100000
                ;mem[2106] <= 30'b000000000000000001010010110000
                ;mem[2107] <= 30'b000000000000000001010011000000
                ;mem[2108] <= 30'b000000000000000001011001000000
                ;mem[2109] <= 30'b000000000000000001011001010000
                ;mem[2110] <= 30'b000000000000000001011001100000
                ;mem[2111] <= 30'b000000000000000001100000000000
                ;mem[2112] <= 30'b000000000000000001100000010000
                ;mem[2113] <= 30'b000000000000000000011111010000
                ;mem[2114] <= 30'b000000000000000000011111100000
                ;mem[2115] <= 30'b000000000000000000011111110000
                ;mem[2116] <= 30'b000000000000000000100000000000
                ;mem[2117] <= 30'b000000000000000000100000010000
                ;mem[2118] <= 30'b000000000000000000100000100000
                ;mem[2119] <= 30'b000000000000000000100000110000
                ;mem[2120] <= 30'b000000000000000000100101010000
                ;mem[2121] <= 30'b000000000000000000100101100000
                ;mem[2122] <= 30'b000000000000000000100101110000
                ;mem[2123] <= 30'b000000000000000000100110000000
                ;mem[2124] <= 30'b000000000000000000100110010000
                ;mem[2125] <= 30'b000000000000000000100110100000
                ;mem[2126] <= 30'b000000000000000000100110110000
                ;mem[2127] <= 30'b000000000000000000100111000000
                ;mem[2128] <= 30'b000000000000000000101100000000
                ;mem[2129] <= 30'b000000000000000000101100010000
                ;mem[2130] <= 30'b000000000000000000101100100000
                ;mem[2131] <= 30'b000000000000000000101100110000
                ;mem[2132] <= 30'b000000000000000000101101000000
                ;mem[2133] <= 30'b000000000000000000110011000000
                ;mem[2134] <= 30'b000000000000000000110011010000
                ;mem[2135] <= 30'b000000000000000000110011100000
                ;mem[2136] <= 30'b000000000000000000111010010000
                ;mem[2137] <= 30'b000000000000000000111010100000
                ;mem[2138] <= 30'b000000001000000000000000000000
                ;mem[2139] <= 30'b000000001000000000000000010000
                ;mem[2140] <= 30'b000000001000000000000000100000
                ;mem[2141] <= 30'b000000001000000000000000110000
                ;mem[2142] <= 30'b000000001000000000000001000000
                ;mem[2143] <= 30'b000000001000000000000111000000
                ;mem[2144] <= 30'b000000001000000000000111010000
                ;mem[2145] <= 30'b000000001000000000000111100000
                ;mem[2146] <= 30'b000000001000000000001110010000
                ;mem[2147] <= 30'b000000001000000000001110100000
                ;mem[2148] <= 30'b000000001000000000010101100000
                ;mem[2149] <= 30'b000000001000000000011100100000
                ;mem[2150] <= 30'b000000001000000000100011010000
                ;mem[2151] <= 30'b000000001000000000100011100000
                ;mem[2152] <= 30'b000000001000000000100011110000
                ;mem[2153] <= 30'b000000001000000000100100000000
                ;mem[2154] <= 30'b000000001000000000100100010000
                ;mem[2155] <= 30'b000000001000000000100100100000
                ;mem[2156] <= 30'b000000001000000000100100110000
                ;mem[2157] <= 30'b000000001000000000101010000000
                ;mem[2158] <= 30'b000000001000000000101010010000
                ;mem[2159] <= 30'b000000001000000000101010100000
                ;mem[2160] <= 30'b000000001000000000101010110000
                ;mem[2161] <= 30'b000000001000000000101011100000
                ;mem[2162] <= 30'b000000001000000000101011110000
                ;mem[2163] <= 30'b000000001000000000101100000000
                ;mem[2164] <= 30'b000000001000000000101100010000
                ;mem[2165] <= 30'b000000001000000000110001000000
                ;mem[2166] <= 30'b000000001000000000110001010000
                ;mem[2167] <= 30'b000000001000000000110011010000
                ;mem[2168] <= 30'b000000001000000000110011100000
                ;mem[2169] <= 30'b000000001000000000110011110000
                ;mem[2170] <= 30'b000000001000000000111010110000
                ;mem[2171] <= 30'b000000001000000000111011000000
                ;mem[2172] <= 30'b000000010000000000000000000000
                ;mem[2173] <= 30'b000000010000000000000000010000
                ;mem[2174] <= 30'b000000010000000000000101000000
                ;mem[2175] <= 30'b000000010000000000000101010000
                ;mem[2176] <= 30'b000000010000000000000111010000
                ;mem[2177] <= 30'b000000010000000000000111100000
                ;mem[2178] <= 30'b000000010000000000000111110000
                ;mem[2179] <= 30'b000000010000000000001110110000
                ;mem[2180] <= 30'b000000010000000000001111000000
                ;mem[2181] <= 30'b000000010000000000010110000000
                ;mem[2182] <= 30'b000000010000000000010110010000
                ;mem[2183] <= 30'b000000010000000000011101010000
                ;mem[2184] <= 30'b000000010000000000011101100000
                ;mem[2185] <= 30'b000000010000000000100100100000
                ;mem[2186] <= 30'b000000010000000000100100110000
                ;mem[2187] <= 30'b000000010000000000101011100000
                ;mem[2188] <= 30'b000000010000000000101011110000
                ;mem[2189] <= 30'b000000010000000000110010100000
                ;mem[2190] <= 30'b000000010000000000110010110000
                ;mem[2191] <= 30'b000000010000000000111001010000
                ;mem[2192] <= 30'b000000010000000000111001100000
                ;mem[2193] <= 30'b000000010000000000111101000000
                ;mem[2194] <= 30'b000000010000000000111101010000
                ;mem[2195] <= 30'b000000010000000000111111110000
                ;mem[2196] <= 30'b000000000000000001000110100000
                ;mem[2197] <= 30'b000000000000000001000110110000
                ;mem[2198] <= 30'b000000000000000001001101010000
                ;mem[2199] <= 30'b000000000000000001001101100000
                ;mem[2200] <= 30'b000000000000000001010001000000
                ;mem[2201] <= 30'b000000000000000001010001010000
                ;mem[2202] <= 30'b000000000000000001010011110000
                ;mem[2203] <= 30'b000000000000000001010100000000
                ;mem[2204] <= 30'b000000000000000001010100010000
                ;mem[2205] <= 30'b000000000000000001011000000000
                ;mem[2206] <= 30'b000000000000000001011000010000
                ;mem[2207] <= 30'b000000000000000001011000100000
                ;mem[2208] <= 30'b000000000000000001011000110000
                ;mem[2209] <= 30'b000000000000000001011001000000
                ;mem[2210] <= 30'b000000000000000001011001010000
                ;mem[2211] <= 30'b000000000000000001011001100000
                ;mem[2212] <= 30'b000000000000000001011001110000
                ;mem[2213] <= 30'b000000000000000001011010000000
                ;mem[2214] <= 30'b000000000000000001011010010000
                ;mem[2215] <= 30'b000000000000000001011010100000
                ;mem[2216] <= 30'b000000000000000001011010110000
                ;mem[2217] <= 30'b000000000000000001011011000000
                ;mem[2218] <= 30'b000000000000000001011111010000
                ;mem[2219] <= 30'b000000000000000001011111100000
                ;mem[2220] <= 30'b000000000000000001011111110000
                ;mem[2221] <= 30'b000000000000000001100000000000
                ;mem[2222] <= 30'b000000000000000001100000010000
                ;mem[2223] <= 30'b000000000000000001100000100000
                ;mem[2224] <= 30'b000000000000000001100000110000
                ;mem[2225] <= 30'b000000000000000001100001000000
                ;mem[2226] <= 30'b000000000000000000101101000000
                ;mem[2227] <= 30'b000000000000000000101101010000
                ;mem[2228] <= 30'b000000000000000000101101100000
                ;mem[2229] <= 30'b000000000000000000101101110000
                ;mem[2230] <= 30'b000000000000000000110011100000
                ;mem[2231] <= 30'b000000000000000000110011110000
                ;mem[2232] <= 30'b000000000000000000110100000000
                ;mem[2233] <= 30'b000000000000000000110100010000
                ;mem[2234] <= 30'b000000000000000000110100100000
                ;mem[2235] <= 30'b000000000000000000110100110000
                ;mem[2236] <= 30'b000000000000000000110101000000
                ;mem[2237] <= 30'b000000000000000000111010010000
                ;mem[2238] <= 30'b000000000000000000111010100000
                ;mem[2239] <= 30'b000000000000000000111010110000
                ;mem[2240] <= 30'b000000000000000000111100000000
                ;mem[2241] <= 30'b000000000000000000111100010000
                ;mem[2242] <= 30'b000000001000000000000001000000
                ;mem[2243] <= 30'b000000001000000000000001010000
                ;mem[2244] <= 30'b000000001000000000000001100000
                ;mem[2245] <= 30'b000000001000000000000001110000
                ;mem[2246] <= 30'b000000001000000000000111100000
                ;mem[2247] <= 30'b000000001000000000000111110000
                ;mem[2248] <= 30'b000000001000000000001000000000
                ;mem[2249] <= 30'b000000001000000000001000010000
                ;mem[2250] <= 30'b000000001000000000001000100000
                ;mem[2251] <= 30'b000000001000000000001000110000
                ;mem[2252] <= 30'b000000001000000000001001000000
                ;mem[2253] <= 30'b000000001000000000001110010000
                ;mem[2254] <= 30'b000000001000000000001110100000
                ;mem[2255] <= 30'b000000001000000000001110110000
                ;mem[2256] <= 30'b000000001000000000010000000000
                ;mem[2257] <= 30'b000000001000000000010000010000
                ;mem[2258] <= 30'b000000001000000000010101000000
                ;mem[2259] <= 30'b000000001000000000010101010000
                ;mem[2260] <= 30'b000000001000000000010101100000
                ;mem[2261] <= 30'b000000001000000000010111110000
                ;mem[2262] <= 30'b000000001000000000011000000000
                ;mem[2263] <= 30'b000000001000000000011100000000
                ;mem[2264] <= 30'b000000001000000000011100010000
                ;mem[2265] <= 30'b000000001000000000011110100000
                ;mem[2266] <= 30'b000000001000000000011110110000
                ;mem[2267] <= 30'b000000001000000000011111000000
                ;mem[2268] <= 30'b000000001000000000100010110000
                ;mem[2269] <= 30'b000000001000000000100011000000
                ;mem[2270] <= 30'b000000001000000000100011010000
                ;mem[2271] <= 30'b000000001000000000100101100000
                ;mem[2272] <= 30'b000000001000000000100101110000
                ;mem[2273] <= 30'b000000001000000000100110000000
                ;mem[2274] <= 30'b000000001000000000101001110000
                ;mem[2275] <= 30'b000000001000000000101010000000
                ;mem[2276] <= 30'b000000001000000000101100100000
                ;mem[2277] <= 30'b000000001000000000101100110000
                ;mem[2278] <= 30'b000000001000000000110000110000
                ;mem[2279] <= 30'b000000001000000000110001000000
                ;mem[2280] <= 30'b000000001000000000110011010000
                ;mem[2281] <= 30'b000000001000000000110011100000
                ;mem[2282] <= 30'b000000001000000000110011110000
                ;mem[2283] <= 30'b000000001000000000110111110000
                ;mem[2284] <= 30'b000000001000000000111000000000
                ;mem[2285] <= 30'b000000001000000000111010010000
                ;mem[2286] <= 30'b000000001000000000111010100000
                ;mem[2287] <= 30'b000000001000000000111010110000
                ;mem[2288] <= 30'b000000001000000000111110110000
                ;mem[2289] <= 30'b000000001000000000111111000000
                ;mem[2290] <= 30'b000000010000000000000000100000
                ;mem[2291] <= 30'b000000010000000000000000110000
                ;mem[2292] <= 30'b000000010000000000000100110000
                ;mem[2293] <= 30'b000000010000000000000101000000
                ;mem[2294] <= 30'b000000010000000000000111010000
                ;mem[2295] <= 30'b000000010000000000000111100000
                ;mem[2296] <= 30'b000000010000000000000111110000
                ;mem[2297] <= 30'b000000010000000000001011110000
                ;mem[2298] <= 30'b000000010000000000001100000000
                ;mem[2299] <= 30'b000000010000000000001110010000
                ;mem[2300] <= 30'b000000010000000000001110100000
                ;mem[2301] <= 30'b000000010000000000001110110000
                ;mem[2302] <= 30'b000000010000000000010010110000
                ;mem[2303] <= 30'b000000010000000000010011000000
                ;mem[2304] <= 30'b000000010000000000010101000000
                ;mem[2305] <= 30'b000000010000000000010101010000
                ;mem[2306] <= 30'b000000010000000000010101100000
                ;mem[2307] <= 30'b000000010000000000011010000000
                ;mem[2308] <= 30'b000000010000000000011010010000
                ;mem[2309] <= 30'b000000010000000000011010100000
                ;mem[2310] <= 30'b000000010000000000011011000000
                ;mem[2311] <= 30'b000000010000000000011011010000
                ;mem[2312] <= 30'b000000010000000000011011100000
                ;mem[2313] <= 30'b000000010000000000011011110000
                ;mem[2314] <= 30'b000000010000000000011100000000
                ;mem[2315] <= 30'b000000010000000000011100010000
                ;mem[2316] <= 30'b000000010000000000011100100000
                ;mem[2317] <= 30'b000000010000000000100001010000
                ;mem[2318] <= 30'b000000010000000000100001100000
                ;mem[2319] <= 30'b000000010000000000100001110000
                ;mem[2320] <= 30'b000000010000000000100010000000
                ;mem[2321] <= 30'b000000010000000000100010010000
                ;mem[2322] <= 30'b000000010000000000100010100000
                ;mem[2323] <= 30'b000000010000000000100011000000
                ;mem[2324] <= 30'b000000010000000000100011010000
                ;mem[2325] <= 30'b000000010000000000100011100000
                ;mem[2326] <= 30'b000000010000000000101010000000
                ;mem[2327] <= 30'b000000010000000000101010010000
                ;mem[2328] <= 30'b000000010000000000110001000000
                ;mem[2329] <= 30'b000000010000000000110001010000
                ;mem[2330] <= 30'b000000010000000000110111110000
                ;mem[2331] <= 30'b000000010000000000111000000000
                ;mem[2332] <= 30'b000000010000000000111000010000
                ;mem[2333] <= 30'b000000010000000000111110110000
                ;mem[2334] <= 30'b000000010000000000111111000000
                ;mem[2335] <= 30'b000000010000000000111111010000
                ;mem[2336] <= 30'b000000000000000001000101000000
                ;mem[2337] <= 30'b000000000000000001000101010000
                ;mem[2338] <= 30'b000000000000000001001011110000
                ;mem[2339] <= 30'b000000000000000001001100000000
                ;mem[2340] <= 30'b000000000000000001001100010000
                ;mem[2341] <= 30'b000000000000000001010010110000
                ;mem[2342] <= 30'b000000000000000001010011000000
                ;mem[2343] <= 30'b000000000000000001010011010000
                ;mem[2344] <= 30'b000000000000000001011001110000
                ;mem[2345] <= 30'b000000000000000001011010000000
                ;mem[2346] <= 30'b000000000000000001100000110000
                ;mem[2347] <= 30'b000000000000000001100001000000
                ;mem[2348] <= 30'b000000000000000001100111100000
                ;mem[2349] <= 30'b000000000000000001100111110000
                ;mem[2350] <= 30'b000000000000000001101000000000
                ;mem[2351] <= 30'b000000000000000001101110100000
                ;mem[2352] <= 30'b000000000000000001101110110000
                ;mem[2353] <= 30'b000000000000000001101111000000
                ;mem[2354] <= 30'b000000000000000000110010010000
                ;mem[2355] <= 30'b000000000000000000110010100000
                ;mem[2356] <= 30'b000000000000000000110010110000
                ;mem[2357] <= 30'b000000000000000000110011000000
                ;mem[2358] <= 30'b000000000000000000110011010000
                ;mem[2359] <= 30'b000000000000000000110011100000
                ;mem[2360] <= 30'b000000000000000000110011110000
                ;mem[2361] <= 30'b000000000000000000110100000000
                ;mem[2362] <= 30'b000000000000000000111001010000
                ;mem[2363] <= 30'b000000000000000000111001100000
                ;mem[2364] <= 30'b000000000000000000111001110000
                ;mem[2365] <= 30'b000000000000000000111010000000
                ;mem[2366] <= 30'b000000000000000000111010010000
                ;mem[2367] <= 30'b000000000000000000111010100000
                ;mem[2368] <= 30'b000000000000000000111010110000
                ;mem[2369] <= 30'b000000000000000000111011000000
                ;mem[2370] <= 30'b000000000000000000111011010000
                ;mem[2371] <= 30'b000000000000000000111011100000
                ;mem[2372] <= 30'b000000000000000000111011110000
                ;mem[2373] <= 30'b000000000000000000111100000000
                ;mem[2374] <= 30'b000000001000000000000110010000
                ;mem[2375] <= 30'b000000001000000000000110100000
                ;mem[2376] <= 30'b000000001000000000000110110000
                ;mem[2377] <= 30'b000000001000000000000111000000
                ;mem[2378] <= 30'b000000001000000000000111010000
                ;mem[2379] <= 30'b000000001000000000000111100000
                ;mem[2380] <= 30'b000000001000000000000111110000
                ;mem[2381] <= 30'b000000001000000000001000000000
                ;mem[2382] <= 30'b000000001000000000001101010000
                ;mem[2383] <= 30'b000000001000000000001101100000
                ;mem[2384] <= 30'b000000001000000000001101110000
                ;mem[2385] <= 30'b000000001000000000001110000000
                ;mem[2386] <= 30'b000000001000000000001110010000
                ;mem[2387] <= 30'b000000001000000000001110100000
                ;mem[2388] <= 30'b000000001000000000001110110000
                ;mem[2389] <= 30'b000000001000000000001111000000
                ;mem[2390] <= 30'b000000001000000000001111010000
                ;mem[2391] <= 30'b000000001000000000001111100000
                ;mem[2392] <= 30'b000000001000000000001111110000
                ;mem[2393] <= 30'b000000001000000000010000000000
                ;mem[2394] <= 30'b000000001000000000010100100000
                ;mem[2395] <= 30'b000000001000000000010101100000
                ;mem[2396] <= 30'b000000001000000000010101110000
                ;mem[2397] <= 30'b000000001000000000010110000000
                ;mem[2398] <= 30'b000000001000000000010110010000
                ;mem[2399] <= 30'b000000001000000000010110100000
                ;mem[2400] <= 30'b000000001000000000010110110000
                ;mem[2401] <= 30'b000000001000000000010111000000
                ;mem[2402] <= 30'b000000001000000000010111010000
                ;mem[2403] <= 30'b000000001000000000010111100000
                ;mem[2404] <= 30'b000000001000000000010111110000
                ;mem[2405] <= 30'b000000001000000000011000000000
                ;mem[2406] <= 30'b000000001000000000011110000000
                ;mem[2407] <= 30'b000000001000000000011110010000
                ;mem[2408] <= 30'b000000001000000000011110100000
                ;mem[2409] <= 30'b000000001000000000011110110000
                ;mem[2410] <= 30'b000000001000000000011111000000
                ;mem[2411] <= 30'b000000001000000000100101100000
                ;mem[2412] <= 30'b000000001000000000100101110000
                ;mem[2413] <= 30'b000000001000000000100110000000
                ;mem[2414] <= 30'b000000001000000000100110010000
                ;mem[2415] <= 30'b000000001000000000101100110000
                ;mem[2416] <= 30'b000000001000000000101101000000
                ;mem[2417] <= 30'b000000001000000000110011110000
                ;mem[2418] <= 30'b000000001000000000110100000000
                ;mem[2419] <= 30'b000000001000000000111010100000
                ;mem[2420] <= 30'b000000001000000000111010110000
                ;mem[2421] <= 30'b000000001000000000111011000000
                ;mem[2422] <= 30'b000000010000000000000000110000
                ;mem[2423] <= 30'b000000010000000000000001000000
                ;mem[2424] <= 30'b000000010000000000000111110000
                ;mem[2425] <= 30'b000000010000000000001000000000
                ;mem[2426] <= 30'b000000010000000000001110100000
                ;mem[2427] <= 30'b000000010000000000001110110000
                ;mem[2428] <= 30'b000000010000000000001111000000
                ;mem[2429] <= 30'b000000010000000000010101100000
                ;mem[2430] <= 30'b000000010000000000010101110000
                ;mem[2431] <= 30'b000000010000000000010110000000
                ;mem[2432] <= 30'b000000010000000000011100010000
                ;mem[2433] <= 30'b000000010000000000011100100000
                ;mem[2434] <= 30'b000000010000000000011100110000
                ;mem[2435] <= 30'b000000010000000000100011000000
                ;mem[2436] <= 30'b000000010000000000100011010000
                ;mem[2437] <= 30'b000000010000000000100011100000
                ;mem[2438] <= 30'b000000010000000000101001110000
                ;mem[2439] <= 30'b000000010000000000101010000000
                ;mem[2440] <= 30'b000000010000000000101010010000
                ;mem[2441] <= 30'b000000010000000000101010100000
                ;mem[2442] <= 30'b000000010000000000110000110000
                ;mem[2443] <= 30'b000000010000000000110001000000
                ;mem[2444] <= 30'b000000010000000000110001010000
                ;mem[2445] <= 30'b000000010000000000110111100000
                ;mem[2446] <= 30'b000000010000000000110111110000
                ;mem[2447] <= 30'b000000010000000000111000000000
                ;mem[2448] <= 30'b000000010000000000111110010000
                ;mem[2449] <= 30'b000000010000000000111110100000
                ;mem[2450] <= 30'b000000010000000000111110110000
                ;mem[2451] <= 30'b000000010000000000111111000000
                ;mem[2452] <= 30'b000000000000000001000100110000
                ;mem[2453] <= 30'b000000000000000001000101000000
                ;mem[2454] <= 30'b000000000000000001000101010000
                ;mem[2455] <= 30'b000000000000000001001011100000
                ;mem[2456] <= 30'b000000000000000001001011110000
                ;mem[2457] <= 30'b000000000000000001001100000000
                ;mem[2458] <= 30'b000000000000000001010010010000
                ;mem[2459] <= 30'b000000000000000001010010100000
                ;mem[2460] <= 30'b000000000000000001010010110000
                ;mem[2461] <= 30'b000000000000000001010011000000
                ;mem[2462] <= 30'b000000000000000001011001010000
                ;mem[2463] <= 30'b000000000000000001011001100000
                ;mem[2464] <= 30'b000000000000000001011001110000
                ;mem[2465] <= 30'b000000000000000001100000000000
                ;mem[2466] <= 30'b000000000000000001100000010000
                ;mem[2467] <= 30'b000000000000000001100000100000
                ;mem[2468] <= 30'b000000000000000001100110110000
                ;mem[2469] <= 30'b000000000000000001100111000000
                ;mem[2470] <= 30'b000000000000000001100111010000
                ;mem[2471] <= 30'b000000000000000001100111100000
                ;mem[2472] <= 30'b000000000000000001101101110000
                ;mem[2473] <= 30'b000000000000000001101110000000
                ;mem[2474] <= 30'b000000000000000001101110010000
                ;mem[2475] <= 30'b000000000000000001110100110000
                ;mem[2476] <= 30'b000000000000000001110101000000
                ;mem[2477] <= 30'b000000000000000000011110000000
                ;mem[2478] <= 30'b000000000000000000011110010000
                ;mem[2479] <= 30'b000000000000000000100100100000
                ;mem[2480] <= 30'b000000000000000000100100110000
                ;mem[2481] <= 30'b000000000000000000100101000000
                ;mem[2482] <= 30'b000000000000000000100101010000
                ;mem[2483] <= 30'b000000000000000000100101100000
                ;mem[2484] <= 30'b000000000000000000100101110000
                ;mem[2485] <= 30'b000000000000000000101011010000
                ;mem[2486] <= 30'b000000000000000000101011100000
                ;mem[2487] <= 30'b000000000000000000101011110000
                ;mem[2488] <= 30'b000000000000000000101100000000
                ;mem[2489] <= 30'b000000000000000000101100010000
                ;mem[2490] <= 30'b000000000000000000101100100000
                ;mem[2491] <= 30'b000000000000000000101100110000
                ;mem[2492] <= 30'b000000000000000000101101000000
                ;mem[2493] <= 30'b000000000000000000110010100000
                ;mem[2494] <= 30'b000000000000000000110010110000
                ;mem[2495] <= 30'b000000000000000000110011000000
                ;mem[2496] <= 30'b000000000000000000110011110000
                ;mem[2497] <= 30'b000000000000000000110100000000
                ;mem[2498] <= 30'b000000000000000000110100010000
                ;mem[2499] <= 30'b000000000000000000110100100000
                ;mem[2500] <= 30'b000000000000000000111001010000
                ;mem[2501] <= 30'b000000000000000000111001100000
                ;mem[2502] <= 30'b000000000000000000111001110000
                ;mem[2503] <= 30'b000000000000000000111011000000
                ;mem[2504] <= 30'b000000000000000000111011010000
                ;mem[2505] <= 30'b000000000000000000111011100000
                ;mem[2506] <= 30'b000000000000000000111011110000
                ;mem[2507] <= 30'b000000001000000000000000000000
                ;mem[2508] <= 30'b000000001000000000000000010000
                ;mem[2509] <= 30'b000000001000000000000000100000
                ;mem[2510] <= 30'b000000001000000000000000110000
                ;mem[2511] <= 30'b000000001000000000000001000000
                ;mem[2512] <= 30'b000000001000000000000110100000
                ;mem[2513] <= 30'b000000001000000000000110110000
                ;mem[2514] <= 30'b000000001000000000000111000000
                ;mem[2515] <= 30'b000000001000000000000111110000
                ;mem[2516] <= 30'b000000001000000000001000000000
                ;mem[2517] <= 30'b000000001000000000001000010000
                ;mem[2518] <= 30'b000000001000000000001000100000
                ;mem[2519] <= 30'b000000001000000000001101010000
                ;mem[2520] <= 30'b000000001000000000001101100000
                ;mem[2521] <= 30'b000000001000000000001101110000
                ;mem[2522] <= 30'b000000001000000000001111000000
                ;mem[2523] <= 30'b000000001000000000001111010000
                ;mem[2524] <= 30'b000000001000000000001111100000
                ;mem[2525] <= 30'b000000001000000000001111110000
                ;mem[2526] <= 30'b000000001000000000010100010000
                ;mem[2527] <= 30'b000000001000000000010100100000
                ;mem[2528] <= 30'b000000001000000000010110010000
                ;mem[2529] <= 30'b000000001000000000010110100000
                ;mem[2530] <= 30'b000000001000000000010110110000
                ;mem[2531] <= 30'b000000001000000000010111000000
                ;mem[2532] <= 30'b000000001000000000011011010000
                ;mem[2533] <= 30'b000000001000000000011011100000
                ;mem[2534] <= 30'b000000001000000000011101100000
                ;mem[2535] <= 30'b000000001000000000011101110000
                ;mem[2536] <= 30'b000000001000000000011110000000
                ;mem[2537] <= 30'b000000001000000000100010010000
                ;mem[2538] <= 30'b000000001000000000100010100000
                ;mem[2539] <= 30'b000000001000000000100011100000
                ;mem[2540] <= 30'b000000001000000000100100100000
                ;mem[2541] <= 30'b000000001000000000100100110000
                ;mem[2542] <= 30'b000000001000000000100101000000
                ;mem[2543] <= 30'b000000001000000000101001100000
                ;mem[2544] <= 30'b000000001000000000101010010000
                ;mem[2545] <= 30'b000000001000000000101010100000
                ;mem[2546] <= 30'b000000001000000000101010110000
                ;mem[2547] <= 30'b000000001000000000101011000000
                ;mem[2548] <= 30'b000000001000000000101011010000
                ;mem[2549] <= 30'b000000001000000000101011100000
                ;mem[2550] <= 30'b000000001000000000101011110000
                ;mem[2551] <= 30'b000000001000000000101100000000
                ;mem[2552] <= 30'b000000001000000000101100010000
                ;mem[2553] <= 30'b000000001000000000110001010000
                ;mem[2554] <= 30'b000000001000000000110001100000
                ;mem[2555] <= 30'b000000001000000000110001110000
                ;mem[2556] <= 30'b000000001000000000110010000000
                ;mem[2557] <= 30'b000000001000000000110010010000
                ;mem[2558] <= 30'b000000001000000000110010100000
                ;mem[2559] <= 30'b000000001000000000110010110000
                ;mem[2560] <= 30'b000000001000000000110011000000
                ;mem[2561] <= 30'b000000001000000000110011010000
                ;mem[2562] <= 30'b000000001000000000110011100000
                ;mem[2563] <= 30'b000000001000000000110011110000
                ;mem[2564] <= 30'b000000001000000000111000100000
                ;mem[2565] <= 30'b000000001000000000111000110000
                ;mem[2566] <= 30'b000000001000000000111001000000
                ;mem[2567] <= 30'b000000001000000000111001010000
                ;mem[2568] <= 30'b000000001000000000111001100000
                ;mem[2569] <= 30'b000000001000000000111001110000
                ;mem[2570] <= 30'b000000001000000000111010000000
                ;mem[2571] <= 30'b000000001000000000111010010000
                ;mem[2572] <= 30'b000000001000000000111010100000
                ;mem[2573] <= 30'b000000001000000000111010110000
                ;mem[2574] <= 30'b000000001000000000111011000000
                ;mem[2575] <= 30'b000000001000000000111011010000
                ;mem[2576] <= 30'b000000010000000000000000000000
                ;mem[2577] <= 30'b000000010000000000000000010000
                ;mem[2578] <= 30'b000000010000000000000101010000
                ;mem[2579] <= 30'b000000010000000000000101100000
                ;mem[2580] <= 30'b000000010000000000000101110000
                ;mem[2581] <= 30'b000000010000000000000110000000
                ;mem[2582] <= 30'b000000010000000000000110010000
                ;mem[2583] <= 30'b000000010000000000000110100000
                ;mem[2584] <= 30'b000000010000000000000110110000
                ;mem[2585] <= 30'b000000010000000000000111000000
                ;mem[2586] <= 30'b000000010000000000000111010000
                ;mem[2587] <= 30'b000000010000000000000111100000
                ;mem[2588] <= 30'b000000010000000000000111110000
                ;mem[2589] <= 30'b000000010000000000001100100000
                ;mem[2590] <= 30'b000000010000000000001100110000
                ;mem[2591] <= 30'b000000010000000000001101000000
                ;mem[2592] <= 30'b000000010000000000001101010000
                ;mem[2593] <= 30'b000000010000000000001101100000
                ;mem[2594] <= 30'b000000010000000000001101110000
                ;mem[2595] <= 30'b000000010000000000001110000000
                ;mem[2596] <= 30'b000000010000000000001110010000
                ;mem[2597] <= 30'b000000010000000000001110100000
                ;mem[2598] <= 30'b000000010000000000001110110000
                ;mem[2599] <= 30'b000000010000000000001111000000
                ;mem[2600] <= 30'b000000010000000000001111010000
                ;mem[2601] <= 30'b000000010000000000010101100000
                ;mem[2602] <= 30'b000000010000000000010101110000
                ;mem[2603] <= 30'b000000010000000000010110000000
                ;mem[2604] <= 30'b000000010000000000010110010000
                ;mem[2605] <= 30'b000000010000000000010110100000
                ;mem[2606] <= 30'b000000010000000000011101000000
                ;mem[2607] <= 30'b000000010000000000011101010000
                ;mem[2608] <= 30'b000000010000000000011101100000
                ;mem[2609] <= 30'b000000010000000000011101110000
                ;mem[2610] <= 30'b000000010000000000100001010000
                ;mem[2611] <= 30'b000000010000000000100001100000
                ;mem[2612] <= 30'b000000010000000000100100010000
                ;mem[2613] <= 30'b000000010000000000100100100000
                ;mem[2614] <= 30'b000000010000000000100100110000
                ;mem[2615] <= 30'b000000010000000000101000010000
                ;mem[2616] <= 30'b000000010000000000101000100000
                ;mem[2617] <= 30'b000000010000000000101000110000
                ;mem[2618] <= 30'b000000010000000000101011100000
                ;mem[2619] <= 30'b000000010000000000101011110000
                ;mem[2620] <= 30'b000000010000000000101100000000
                ;mem[2621] <= 30'b000000010000000000101111100000
                ;mem[2622] <= 30'b000000010000000000101111110000
                ;mem[2623] <= 30'b000000010000000000110010100000
                ;mem[2624] <= 30'b000000010000000000110010110000
                ;mem[2625] <= 30'b000000010000000000110011000000
                ;mem[2626] <= 30'b000000010000000000110110100000
                ;mem[2627] <= 30'b000000010000000000110110110000
                ;mem[2628] <= 30'b000000010000000000110111000000
                ;mem[2629] <= 30'b000000010000000000110111010000
                ;mem[2630] <= 30'b000000010000000000111001000000
                ;mem[2631] <= 30'b000000010000000000111001010000
                ;mem[2632] <= 30'b000000010000000000111001100000
                ;mem[2633] <= 30'b000000010000000000111001110000
                ;mem[2634] <= 30'b000000010000000000111010000000
                ;mem[2635] <= 30'b000000010000000000111101110000
                ;mem[2636] <= 30'b000000010000000000111110000000
                ;mem[2637] <= 30'b000000010000000000111110010000
                ;mem[2638] <= 30'b000000010000000000111110100000
                ;mem[2639] <= 30'b000000010000000000111110110000
                ;mem[2640] <= 30'b000000010000000000111111000000
                ;mem[2641] <= 30'b000000010000000000111111010000
                ;mem[2642] <= 30'b000000010000000000111111100000
                ;mem[2643] <= 30'b000000010000000000111111110000
                ;mem[2644] <= 30'b000000000000000001000000000000
                ;mem[2645] <= 30'b000000000000000001000011100000
                ;mem[2646] <= 30'b000000000000000001000011110000
                ;mem[2647] <= 30'b000000000000000001000110100000
                ;mem[2648] <= 30'b000000000000000001000110110000
                ;mem[2649] <= 30'b000000000000000001000111000000
                ;mem[2650] <= 30'b000000000000000001001010100000
                ;mem[2651] <= 30'b000000000000000001001010110000
                ;mem[2652] <= 30'b000000000000000001001011000000
                ;mem[2653] <= 30'b000000000000000001001011010000
                ;mem[2654] <= 30'b000000000000000001001101000000
                ;mem[2655] <= 30'b000000000000000001001101010000
                ;mem[2656] <= 30'b000000000000000001001101100000
                ;mem[2657] <= 30'b000000000000000001001101110000
                ;mem[2658] <= 30'b000000000000000001001110000000
                ;mem[2659] <= 30'b000000000000000001010001110000
                ;mem[2660] <= 30'b000000000000000001010010000000
                ;mem[2661] <= 30'b000000000000000001010010010000
                ;mem[2662] <= 30'b000000000000000001010010100000
                ;mem[2663] <= 30'b000000000000000001010010110000
                ;mem[2664] <= 30'b000000000000000001010011000000
                ;mem[2665] <= 30'b000000000000000001010011010000
                ;mem[2666] <= 30'b000000000000000001010011100000
                ;mem[2667] <= 30'b000000000000000001010011110000
                ;mem[2668] <= 30'b000000000000000001010100000000
                ;mem[2669] <= 30'b000000000000000001010100010000
                ;mem[2670] <= 30'b000000000000000001010100100000
                ;mem[2671] <= 30'b000000000000000001010100110000
                ;mem[2672] <= 30'b000000000000000001011001010000
                ;mem[2673] <= 30'b000000000000000001011001100000
                ;mem[2674] <= 30'b000000000000000001011001110000
                ;mem[2675] <= 30'b000000000000000001011010000000
                ;mem[2676] <= 30'b000000000000000001011010010000
                ;mem[2677] <= 30'b000000000000000001011010100000
                ;mem[2678] <= 30'b000000000000000001011010110000
                ;mem[2679] <= 30'b000000000000000001011011000000
                ;mem[2680] <= 30'b000000000000000001011011010000
                ;mem[2681] <= 30'b000000000000000001100001000000
                ;mem[2682] <= 30'b000000000000000000100111100000
                ;mem[2683] <= 30'b000000000000000000101110100000
                ;mem[2684] <= 30'b000000000000000000110101100000
                ;mem[2685] <= 30'b000000000000000000111010100000
                ;mem[2686] <= 30'b000000000000000000111100100000
                ;mem[2687] <= 30'b000000001000000000000010100000
                ;mem[2688] <= 30'b000000001000000000001001100000
                ;mem[2689] <= 30'b000000001000000000001110100000
                ;mem[2690] <= 30'b000000001000000000010000100000
                ;mem[2691] <= 30'b000000001000000000010101100000
                ;mem[2692] <= 30'b000000001000000000010111100000
                ;mem[2693] <= 30'b000000001000000000011100010000
                ;mem[2694] <= 30'b000000001000000000011100100000
                ;mem[2695] <= 30'b000000001000000000011110010000
                ;mem[2696] <= 30'b000000001000000000011110100000
                ;mem[2697] <= 30'b000000001000000000100011010000
                ;mem[2698] <= 30'b000000001000000000100011100000
                ;mem[2699] <= 30'b000000001000000000100101010000
                ;mem[2700] <= 30'b000000001000000000100101100000
                ;mem[2701] <= 30'b000000001000000000101010010000
                ;mem[2702] <= 30'b000000001000000000101100010000
                ;mem[2703] <= 30'b000000001000000000101100100000
                ;mem[2704] <= 30'b000000001000000000110001010000
                ;mem[2705] <= 30'b000000001000000000110011010000
                ;mem[2706] <= 30'b000000001000000000111000000000
                ;mem[2707] <= 30'b000000001000000000111000010000
                ;mem[2708] <= 30'b000000001000000000111000110000
                ;mem[2709] <= 30'b000000001000000000111001000000
                ;mem[2710] <= 30'b000000001000000000111001010000
                ;mem[2711] <= 30'b000000001000000000111001100000
                ;mem[2712] <= 30'b000000001000000000111001110000
                ;mem[2713] <= 30'b000000001000000000111010000000
                ;mem[2714] <= 30'b000000001000000000111010010000
                ;mem[2715] <= 30'b000000001000000000111111000000
                ;mem[2716] <= 30'b000000001000000000111111010000
                ;mem[2717] <= 30'b000000001000000000111111100000
                ;mem[2718] <= 30'b000000001000000000111111110000
                ;mem[2719] <= 30'b000000010000000000000000010000
                ;mem[2720] <= 30'b000000010000000000000000100000
                ;mem[2721] <= 30'b000000010000000000000101010000
                ;mem[2722] <= 30'b000000010000000000000111010000
                ;mem[2723] <= 30'b000000010000000000001100000000
                ;mem[2724] <= 30'b000000010000000000001100010000
                ;mem[2725] <= 30'b000000010000000000001100110000
                ;mem[2726] <= 30'b000000010000000000001101000000
                ;mem[2727] <= 30'b000000010000000000001101010000
                ;mem[2728] <= 30'b000000010000000000001101100000
                ;mem[2729] <= 30'b000000010000000000001101110000
                ;mem[2730] <= 30'b000000010000000000001110000000
                ;mem[2731] <= 30'b000000010000000000001110010000
                ;mem[2732] <= 30'b000000010000000000010011000000
                ;mem[2733] <= 30'b000000010000000000010011010000
                ;mem[2734] <= 30'b000000010000000000010011100000
                ;mem[2735] <= 30'b000000010000000000010011110000
                ;mem[2736] <= 30'b000000010000000000010100000000
                ;mem[2737] <= 30'b000000010000000000010100010000
                ;mem[2738] <= 30'b000000010000000000010100100000
                ;mem[2739] <= 30'b000000010000000000010100110000
                ;mem[2740] <= 30'b000000010000000000010101000000
                ;mem[2741] <= 30'b000000010000000000010101010000
                ;mem[2742] <= 30'b000000010000000000010101100000
                ;mem[2743] <= 30'b000000010000000000011010000000
                ;mem[2744] <= 30'b000000010000000000011010010000
                ;mem[2745] <= 30'b000000010000000000011100000000
                ;mem[2746] <= 30'b000000010000000000011100010000
                ;mem[2747] <= 30'b000000010000000000011100100000
                ;mem[2748] <= 30'b000000010000000000011100110000
                ;mem[2749] <= 30'b000000010000000000100011000000
                ;mem[2750] <= 30'b000000010000000000100011010000
                ;mem[2751] <= 30'b000000010000000000101010000000
                ;mem[2752] <= 30'b000000010000000000101010010000
                ;mem[2753] <= 30'b000000010000000000110001000000
                ;mem[2754] <= 30'b000000010000000000111000000000
                ;mem[2755] <= 30'b000000010000000000111111000000
                ;mem[2756] <= 30'b000000000000000001000101000000
                ;mem[2757] <= 30'b000000000000000001001100000000
                ;mem[2758] <= 30'b000000000000000001010011000000
                ;mem[2759] <= 30'b000000000000000001011001110000
                ;mem[2760] <= 30'b000000000000000001011010000000
                ;mem[2761] <= 30'b000000000000000001100000110000
                ;mem[2762] <= 30'b000000000000000001100001000000
                ;mem[2763] <= 30'b000000000000000001101000000000
                ;mem[2764] <= 30'b000000000000000000101110000000
                ;mem[2765] <= 30'b000000000000000000101110010000
                ;mem[2766] <= 30'b000000000000000000110100100000
                ;mem[2767] <= 30'b000000000000000000110100110000
                ;mem[2768] <= 30'b000000000000000000110101000000
                ;mem[2769] <= 30'b000000000000000000110101010000
                ;mem[2770] <= 30'b000000000000000000110101100000
                ;mem[2771] <= 30'b000000000000000000111011010000
                ;mem[2772] <= 30'b000000000000000000111011100000
                ;mem[2773] <= 30'b000000000000000000111011110000
                ;mem[2774] <= 30'b000000000000000000111100000000
                ;mem[2775] <= 30'b000000000000000000111100010000
                ;mem[2776] <= 30'b000000000000000000111100100000
                ;mem[2777] <= 30'b000000000000000000111100110000
                ;mem[2778] <= 30'b000000000000000000111101000000
                ;mem[2779] <= 30'b000000000000000000111101010000
                ;mem[2780] <= 30'b000000001000000000000010000000
                ;mem[2781] <= 30'b000000001000000000000010010000
                ;mem[2782] <= 30'b000000001000000000001000100000
                ;mem[2783] <= 30'b000000001000000000001000110000
                ;mem[2784] <= 30'b000000001000000000001001000000
                ;mem[2785] <= 30'b000000001000000000001001010000
                ;mem[2786] <= 30'b000000001000000000001001100000
                ;mem[2787] <= 30'b000000001000000000001111010000
                ;mem[2788] <= 30'b000000001000000000001111100000
                ;mem[2789] <= 30'b000000001000000000001111110000
                ;mem[2790] <= 30'b000000001000000000010000000000
                ;mem[2791] <= 30'b000000001000000000010000010000
                ;mem[2792] <= 30'b000000001000000000010000100000
                ;mem[2793] <= 30'b000000001000000000010000110000
                ;mem[2794] <= 30'b000000001000000000010001000000
                ;mem[2795] <= 30'b000000001000000000010001010000
                ;mem[2796] <= 30'b000000001000000000010101110000
                ;mem[2797] <= 30'b000000001000000000010110000000
                ;mem[2798] <= 30'b000000001000000000010110010000
                ;mem[2799] <= 30'b000000001000000000010110100000
                ;mem[2800] <= 30'b000000001000000000010110110000
                ;mem[2801] <= 30'b000000001000000000010111000000
                ;mem[2802] <= 30'b000000001000000000010111010000
                ;mem[2803] <= 30'b000000001000000000010111100000
                ;mem[2804] <= 30'b000000001000000000010111110000
                ;mem[2805] <= 30'b000000001000000000011000000000
                ;mem[2806] <= 30'b000000001000000000011000010000
                ;mem[2807] <= 30'b000000001000000000011100100000
                ;mem[2808] <= 30'b000000001000000000011100110000
                ;mem[2809] <= 30'b000000001000000000011101000000
                ;mem[2810] <= 30'b000000001000000000011101010000
                ;mem[2811] <= 30'b000000001000000000011110000000
                ;mem[2812] <= 30'b000000001000000000011110010000
                ;mem[2813] <= 30'b000000001000000000011110100000
                ;mem[2814] <= 30'b000000001000000000011110110000
                ;mem[2815] <= 30'b000000001000000000011111000000
                ;mem[2816] <= 30'b000000001000000000100011010000
                ;mem[2817] <= 30'b000000001000000000100011100000
                ;mem[2818] <= 30'b000000001000000000100011110000
                ;mem[2819] <= 30'b000000001000000000100100000000
                ;mem[2820] <= 30'b000000001000000000100100110000
                ;mem[2821] <= 30'b000000001000000000100101000000
                ;mem[2822] <= 30'b000000001000000000100101010000
                ;mem[2823] <= 30'b000000001000000000100101100000
                ;mem[2824] <= 30'b000000001000000000100101110000
                ;mem[2825] <= 30'b000000001000000000100110000000
                ;mem[2826] <= 30'b000000001000000000101010010000
                ;mem[2827] <= 30'b000000001000000000101010100000
                ;mem[2828] <= 30'b000000001000000000101010110000
                ;mem[2829] <= 30'b000000001000000000101011010000
                ;mem[2830] <= 30'b000000001000000000101011100000
                ;mem[2831] <= 30'b000000001000000000101011110000
                ;mem[2832] <= 30'b000000001000000000101100000000
                ;mem[2833] <= 30'b000000001000000000101100010000
                ;mem[2834] <= 30'b000000001000000000101100100000
                ;mem[2835] <= 30'b000000001000000000101100110000
                ;mem[2836] <= 30'b000000001000000000110001000000
                ;mem[2837] <= 30'b000000001000000000110001010000
                ;mem[2838] <= 30'b000000001000000000110001100000
                ;mem[2839] <= 30'b000000001000000000110001110000
                ;mem[2840] <= 30'b000000001000000000110010000000
                ;mem[2841] <= 30'b000000001000000000110010010000
                ;mem[2842] <= 30'b000000001000000000110010100000
                ;mem[2843] <= 30'b000000001000000000110010110000
                ;mem[2844] <= 30'b000000001000000000110011000000
                ;mem[2845] <= 30'b000000001000000000110011010000
                ;mem[2846] <= 30'b000000001000000000110011100000
                ;mem[2847] <= 30'b000000001000000000111000000000
                ;mem[2848] <= 30'b000000001000000000111000010000
                ;mem[2849] <= 30'b000000001000000000111000100000
                ;mem[2850] <= 30'b000000001000000000111000110000
                ;mem[2851] <= 30'b000000001000000000111001000000
                ;mem[2852] <= 30'b000000001000000000111001010000
                ;mem[2853] <= 30'b000000001000000000111010000000
                ;mem[2854] <= 30'b000000001000000000111010010000
                ;mem[2855] <= 30'b000000001000000000111010100000
                ;mem[2856] <= 30'b000000010000000000000000000000
                ;mem[2857] <= 30'b000000010000000000000000010000
                ;mem[2858] <= 30'b000000010000000000000000100000
                ;mem[2859] <= 30'b000000010000000000000000110000
                ;mem[2860] <= 30'b000000010000000000000101000000
                ;mem[2861] <= 30'b000000010000000000000101010000
                ;mem[2862] <= 30'b000000010000000000000101100000
                ;mem[2863] <= 30'b000000010000000000000101110000
                ;mem[2864] <= 30'b000000010000000000000110000000
                ;mem[2865] <= 30'b000000010000000000000110010000
                ;mem[2866] <= 30'b000000010000000000000110100000
                ;mem[2867] <= 30'b000000010000000000000110110000
                ;mem[2868] <= 30'b000000010000000000000111000000
                ;mem[2869] <= 30'b000000010000000000000111010000
                ;mem[2870] <= 30'b000000010000000000000111100000
                ;mem[2871] <= 30'b000000010000000000001100000000
                ;mem[2872] <= 30'b000000010000000000001100010000
                ;mem[2873] <= 30'b000000010000000000001100100000
                ;mem[2874] <= 30'b000000010000000000001100110000
                ;mem[2875] <= 30'b000000010000000000001101000000
                ;mem[2876] <= 30'b000000010000000000001101010000
                ;mem[2877] <= 30'b000000010000000000001110000000
                ;mem[2878] <= 30'b000000010000000000001110010000
                ;mem[2879] <= 30'b000000010000000000001110100000
                ;mem[2880] <= 30'b000000010000000000010100110000
                ;mem[2881] <= 30'b000000010000000000010101000000
                ;mem[2882] <= 30'b000000010000000000010101010000
                ;mem[2883] <= 30'b000000010000000000011011110000
                ;mem[2884] <= 30'b000000010000000000011100000000
                ;mem[2885] <= 30'b000000010000000000011100010000
                ;mem[2886] <= 30'b000000010000000000100010100000
                ;mem[2887] <= 30'b000000010000000000100010110000
                ;mem[2888] <= 30'b000000010000000000100011000000
                ;mem[2889] <= 30'b000000010000000000101001010000
                ;mem[2890] <= 30'b000000010000000000101001100000
                ;mem[2891] <= 30'b000000010000000000101001110000
                ;mem[2892] <= 30'b000000010000000000110000010000
                ;mem[2893] <= 30'b000000010000000000110000100000
                ;mem[2894] <= 30'b000000010000000000110000110000
                ;mem[2895] <= 30'b000000010000000000110111000000
                ;mem[2896] <= 30'b000000010000000000110111010000
                ;mem[2897] <= 30'b000000010000000000110111100000
                ;mem[2898] <= 30'b000000010000000000111110000000
                ;mem[2899] <= 30'b000000010000000000111110010000
                ;mem[2900] <= 30'b000000000000000001000100010000
                ;mem[2901] <= 30'b000000000000000001000100100000
                ;mem[2902] <= 30'b000000000000000001000100110000
                ;mem[2903] <= 30'b000000000000000001001011000000
                ;mem[2904] <= 30'b000000000000000001001011010000
                ;mem[2905] <= 30'b000000000000000001001011100000
                ;mem[2906] <= 30'b000000000000000001010010000000
                ;mem[2907] <= 30'b000000000000000001010010010000
                ;mem[2908] <= 30'b000000000000000001011000110000
                ;mem[2909] <= 30'b000000000000000001011001000000
                ;mem[2910] <= 30'b000000000000000001011001010000
                ;mem[2911] <= 30'b000000000000000001011111100000
                ;mem[2912] <= 30'b000000000000000001011111110000
                ;mem[2913] <= 30'b000000000000000001100000000000
                ;mem[2914] <= 30'b000000000000000001100000010000
                ;mem[2915] <= 30'b000000000000000001100110100000
                ;mem[2916] <= 30'b000000000000000001100110110000
                ;mem[2917] <= 30'b000000000000000001100111000000
                ;mem[2918] <= 30'b000000000000000001101101100000
                ;mem[2919] <= 30'b000000000000000000011000010000
                ;mem[2920] <= 30'b000000000000000000011000100000
                ;mem[2921] <= 30'b000000000000000000011000110000
                ;mem[2922] <= 30'b000000000000000000011111000000
                ;mem[2923] <= 30'b000000000000000000011111010000
                ;mem[2924] <= 30'b000000000000000000011111100000
                ;mem[2925] <= 30'b000000000000000000011111110000
                ;mem[2926] <= 30'b000000000000000000100000000000
                ;mem[2927] <= 30'b000000000000000000100110000000
                ;mem[2928] <= 30'b000000000000000000100110010000
                ;mem[2929] <= 30'b000000000000000000100110100000
                ;mem[2930] <= 30'b000000000000000000101100110000
                ;mem[2931] <= 30'b000000000000000000101101000000
                ;mem[2932] <= 30'b000000000000000000101101010000
                ;mem[2933] <= 30'b000000000000000000110011110000
                ;mem[2934] <= 30'b000000000000000000110100000000
                ;mem[2935] <= 30'b000000000000000000111010100000
                ;mem[2936] <= 30'b000000000000000000111010110000
                ;mem[2937] <= 30'b000000000000000000111011000000
                ;mem[2938] <= 30'b000000001000000000000000110000
                ;mem[2939] <= 30'b000000001000000000000001000000
                ;mem[2940] <= 30'b000000001000000000000001010000
                ;mem[2941] <= 30'b000000001000000000000111110000
                ;mem[2942] <= 30'b000000001000000000001000000000
                ;mem[2943] <= 30'b000000001000000000001110100000
                ;mem[2944] <= 30'b000000001000000000001110110000
                ;mem[2945] <= 30'b000000001000000000001111000000
                ;mem[2946] <= 30'b000000001000000000010101100000
                ;mem[2947] <= 30'b000000001000000000010101110000
                ;mem[2948] <= 30'b000000001000000000011100100000
                ;mem[2949] <= 30'b000000001000000000011100110000
                ;mem[2950] <= 30'b000000001000000000100011010000
                ;mem[2951] <= 30'b000000001000000000100011100000
                ;mem[2952] <= 30'b000000001000000000100011110000
                ;mem[2953] <= 30'b000000001000000000101010010000
                ;mem[2954] <= 30'b000000001000000000101010100000
                ;mem[2955] <= 30'b000000001000000000110001010000
                ;mem[2956] <= 30'b000000001000000000110001100000
                ;mem[2957] <= 30'b000000001000000000110001110000
                ;mem[2958] <= 30'b000000001000000000110010000000
                ;mem[2959] <= 30'b000000001000000000110010010000
                ;mem[2960] <= 30'b000000001000000000110010100000
                ;mem[2961] <= 30'b000000001000000000110010110000
                ;mem[2962] <= 30'b000000001000000000110011000000
                ;mem[2963] <= 30'b000000001000000000110011010000
                ;mem[2964] <= 30'b000000001000000000111000010000
                ;mem[2965] <= 30'b000000001000000000111000100000
                ;mem[2966] <= 30'b000000001000000000111000110000
                ;mem[2967] <= 30'b000000001000000000111001000000
                ;mem[2968] <= 30'b000000001000000000111001010000
                ;mem[2969] <= 30'b000000001000000000111001100000
                ;mem[2970] <= 30'b000000001000000000111001110000
                ;mem[2971] <= 30'b000000001000000000111010000000
                ;mem[2972] <= 30'b000000001000000000111010010000
                ;mem[2973] <= 30'b000000001000000000111010100000
                ;mem[2974] <= 30'b000000001000000000111111010000
                ;mem[2975] <= 30'b000000001000000000111111100000
                ;mem[2976] <= 30'b000000001000000000111111110000
                ;mem[2977] <= 30'b000000010000000000000101010000
                ;mem[2978] <= 30'b000000010000000000000101100000
                ;mem[2979] <= 30'b000000010000000000000101110000
                ;mem[2980] <= 30'b000000010000000000000110000000
                ;mem[2981] <= 30'b000000010000000000000110010000
                ;mem[2982] <= 30'b000000010000000000000110100000
                ;mem[2983] <= 30'b000000010000000000000110110000
                ;mem[2984] <= 30'b000000010000000000000111000000
                ;mem[2985] <= 30'b000000010000000000000111010000
                ;mem[2986] <= 30'b000000010000000000001100010000
                ;mem[2987] <= 30'b000000010000000000001100100000
                ;mem[2988] <= 30'b000000010000000000001100110000
                ;mem[2989] <= 30'b000000010000000000001101000000
                ;mem[2990] <= 30'b000000010000000000001101010000
                ;mem[2991] <= 30'b000000010000000000001101100000
                ;mem[2992] <= 30'b000000010000000000001101110000
                ;mem[2993] <= 30'b000000010000000000001110000000
                ;mem[2994] <= 30'b000000010000000000001110010000
                ;mem[2995] <= 30'b000000010000000000001110100000
                ;mem[2996] <= 30'b000000010000000000010011010000
                ;mem[2997] <= 30'b000000010000000000010011100000
                ;mem[2998] <= 30'b000000010000000000010011110000
                ;mem[2999] <= 30'b000000010000000000010100000000
                ;mem[3000] <= 30'b000000010000000000010101010000
                ;mem[3001] <= 30'b000000010000000000010101100000
                ;mem[3002] <= 30'b000000010000000000010101110000
                ;mem[3003] <= 30'b000000010000000000011010010000
                ;mem[3004] <= 30'b000000010000000000011010100000
                ;mem[3005] <= 30'b000000010000000000011010110000
                ;mem[3006] <= 30'b000000010000000000011100100000
                ;mem[3007] <= 30'b000000010000000000011100110000
                ;mem[3008] <= 30'b000000010000000000100001100000
                ;mem[3009] <= 30'b000000010000000000100001110000
                ;mem[3010] <= 30'b000000010000000000100011100000
                ;mem[3011] <= 30'b000000010000000000100011110000
                ;mem[3012] <= 30'b000000010000000000101000100000
                ;mem[3013] <= 30'b000000010000000000101000110000
                ;mem[3014] <= 30'b000000010000000000101010100000
                ;mem[3015] <= 30'b000000010000000000101010110000
                ;mem[3016] <= 30'b000000010000000000101111100000
                ;mem[3017] <= 30'b000000010000000000101111110000
                ;mem[3018] <= 30'b000000010000000000110000000000
                ;mem[3019] <= 30'b000000010000000000110001010000
                ;mem[3020] <= 30'b000000010000000000110001100000
                ;mem[3021] <= 30'b000000010000000000110001110000
                ;mem[3022] <= 30'b000000010000000000110110110000
                ;mem[3023] <= 30'b000000010000000000110111000000
                ;mem[3024] <= 30'b000000010000000000110111010000
                ;mem[3025] <= 30'b000000010000000000111000000000
                ;mem[3026] <= 30'b000000010000000000111000010000
                ;mem[3027] <= 30'b000000010000000000111000100000
                ;mem[3028] <= 30'b000000010000000000111000110000
                ;mem[3029] <= 30'b000000010000000000111110000000
                ;mem[3030] <= 30'b000000010000000000111110010000
                ;mem[3031] <= 30'b000000010000000000111110100000
                ;mem[3032] <= 30'b000000010000000000111110110000
                ;mem[3033] <= 30'b000000010000000000111111000000
                ;mem[3034] <= 30'b000000010000000000111111010000
                ;mem[3035] <= 30'b000000000000000001000011100000
                ;mem[3036] <= 30'b000000000000000001000011110000
                ;mem[3037] <= 30'b000000000000000001000100000000
                ;mem[3038] <= 30'b000000000000000001000101010000
                ;mem[3039] <= 30'b000000000000000001000101100000
                ;mem[3040] <= 30'b000000000000000001000101110000
                ;mem[3041] <= 30'b000000000000000001001010110000
                ;mem[3042] <= 30'b000000000000000001001011000000
                ;mem[3043] <= 30'b000000000000000001001011010000
                ;mem[3044] <= 30'b000000000000000001001100000000
                ;mem[3045] <= 30'b000000000000000001001100010000
                ;mem[3046] <= 30'b000000000000000001001100100000
                ;mem[3047] <= 30'b000000000000000001001100110000
                ;mem[3048] <= 30'b000000000000000001010010000000
                ;mem[3049] <= 30'b000000000000000001010010010000
                ;mem[3050] <= 30'b000000000000000001010010100000
                ;mem[3051] <= 30'b000000000000000001010010110000
                ;mem[3052] <= 30'b000000000000000001010011000000
                ;mem[3053] <= 30'b000000000000000001010011010000
                ;mem[3054] <= 30'b000000000000000001011001010000
                ;mem[3055] <= 30'b000000000000000001011001100000
                ;mem[3056] <= 30'b000000000000000001011001110000
                ;mem[3057] <= 30'b000000000000000000010111100000
                ;mem[3058] <= 30'b000000000000000000011110010000
                ;mem[3059] <= 30'b000000000000000000011110100000
                ;mem[3060] <= 30'b000000000000000000100101010000
                ;mem[3061] <= 30'b000000000000000000101100010000
                ;mem[3062] <= 30'b000000000000000000110011000000
                ;mem[3063] <= 30'b000000000000000000110011010000
                ;mem[3064] <= 30'b000000000000000000111010000000
                ;mem[3065] <= 30'b000000000000000000111010010000
                ;mem[3066] <= 30'b000000001000000000000000010000
                ;mem[3067] <= 30'b000000001000000000000111000000
                ;mem[3068] <= 30'b000000001000000000000111010000
                ;mem[3069] <= 30'b000000001000000000001110000000
                ;mem[3070] <= 30'b000000001000000000001110010000
                ;mem[3071] <= 30'b000000001000000000010100110000
                ;mem[3072] <= 30'b000000001000000000010101000000
                ;mem[3073] <= 30'b000000001000000000010101010000
                ;mem[3074] <= 30'b000000001000000000010111110000
                ;mem[3075] <= 30'b000000001000000000011011110000
                ;mem[3076] <= 30'b000000001000000000011100000000
                ;mem[3077] <= 30'b000000001000000000011110000000
                ;mem[3078] <= 30'b000000001000000000011110010000
                ;mem[3079] <= 30'b000000001000000000011110100000
                ;mem[3080] <= 30'b000000001000000000011110110000
                ;mem[3081] <= 30'b000000001000000000011111000000
                ;mem[3082] <= 30'b000000001000000000100010110000
                ;mem[3083] <= 30'b000000001000000000100011000000
                ;mem[3084] <= 30'b000000001000000000100100110000
                ;mem[3085] <= 30'b000000001000000000100101000000
                ;mem[3086] <= 30'b000000001000000000100101010000
                ;mem[3087] <= 30'b000000001000000000100110000000
                ;mem[3088] <= 30'b000000001000000000100110010000
                ;mem[3089] <= 30'b000000001000000000101001110000
                ;mem[3090] <= 30'b000000001000000000101010000000
                ;mem[3091] <= 30'b000000001000000000101011110000
                ;mem[3092] <= 30'b000000001000000000101100000000
                ;mem[3093] <= 30'b000000001000000000101101000000
                ;mem[3094] <= 30'b000000001000000000101101010000
                ;mem[3095] <= 30'b000000001000000000110000110000
                ;mem[3096] <= 30'b000000001000000000110001000000
                ;mem[3097] <= 30'b000000001000000000110010100000
                ;mem[3098] <= 30'b000000001000000000110010110000
                ;mem[3099] <= 30'b000000001000000000110100000000
                ;mem[3100] <= 30'b000000001000000000110100010000
                ;mem[3101] <= 30'b000000001000000000110111110000
                ;mem[3102] <= 30'b000000001000000000111000000000
                ;mem[3103] <= 30'b000000001000000000111001100000
                ;mem[3104] <= 30'b000000001000000000111001110000
                ;mem[3105] <= 30'b000000001000000000111011000000
                ;mem[3106] <= 30'b000000001000000000111011010000
                ;mem[3107] <= 30'b000000001000000000111111000000
                ;mem[3108] <= 30'b000000001000000000111111010000
                ;mem[3109] <= 30'b000000010000000000000000000000
                ;mem[3110] <= 30'b000000010000000000000001000000
                ;mem[3111] <= 30'b000000010000000000000001010000
                ;mem[3112] <= 30'b000000010000000000000100110000
                ;mem[3113] <= 30'b000000010000000000000101000000
                ;mem[3114] <= 30'b000000010000000000000110100000
                ;mem[3115] <= 30'b000000010000000000000110110000
                ;mem[3116] <= 30'b000000010000000000001000000000
                ;mem[3117] <= 30'b000000010000000000001000010000
                ;mem[3118] <= 30'b000000010000000000001011110000
                ;mem[3119] <= 30'b000000010000000000001100000000
                ;mem[3120] <= 30'b000000010000000000001101100000
                ;mem[3121] <= 30'b000000010000000000001101110000
                ;mem[3122] <= 30'b000000010000000000001111000000
                ;mem[3123] <= 30'b000000010000000000001111010000
                ;mem[3124] <= 30'b000000010000000000010011000000
                ;mem[3125] <= 30'b000000010000000000010011010000
                ;mem[3126] <= 30'b000000010000000000010100010000
                ;mem[3127] <= 30'b000000010000000000010100100000
                ;mem[3128] <= 30'b000000010000000000010110000000
                ;mem[3129] <= 30'b000000010000000000010110010000
                ;mem[3130] <= 30'b000000010000000000011010000000
                ;mem[3131] <= 30'b000000010000000000011010010000
                ;mem[3132] <= 30'b000000010000000000011011010000
                ;mem[3133] <= 30'b000000010000000000011011100000
                ;mem[3134] <= 30'b000000010000000000011101000000
                ;mem[3135] <= 30'b000000010000000000100001010000
                ;mem[3136] <= 30'b000000010000000000100001100000
                ;mem[3137] <= 30'b000000010000000000100001110000
                ;mem[3138] <= 30'b000000010000000000100010010000
                ;mem[3139] <= 30'b000000010000000000100010100000
                ;mem[3140] <= 30'b000000010000000000100011110000
                ;mem[3141] <= 30'b000000010000000000100100000000
                ;mem[3142] <= 30'b000000010000000000101000100000
                ;mem[3143] <= 30'b000000010000000000101000110000
                ;mem[3144] <= 30'b000000010000000000101001000000
                ;mem[3145] <= 30'b000000010000000000101001010000
                ;mem[3146] <= 30'b000000010000000000101001100000
                ;mem[3147] <= 30'b000000010000000000101010010000
                ;mem[3148] <= 30'b000000010000000000101010100000
                ;mem[3149] <= 30'b000000010000000000101010110000
                ;mem[3150] <= 30'b000000010000000000101111110000
                ;mem[3151] <= 30'b000000010000000000110000000000
                ;mem[3152] <= 30'b000000010000000000110000010000
                ;mem[3153] <= 30'b000000010000000000110000100000
                ;mem[3154] <= 30'b000000010000000000110000110000
                ;mem[3155] <= 30'b000000010000000000110001000000
                ;mem[3156] <= 30'b000000010000000000110001010000
                ;mem[3157] <= 30'b000000010000000000110001100000
                ;mem[3158] <= 30'b000000010000000000110111010000
                ;mem[3159] <= 30'b000000010000000000110111100000
                ;mem[3160] <= 30'b000000010000000000110111110000
                ;mem[3161] <= 30'b000000010000000000111000000000
                ;mem[3162] <= 30'b000000010000000000111110010000
                ;mem[3163] <= 30'b000000010000000000111110100000
                ;mem[3164] <= 30'b000000010000000000111110110000
                ;mem[3165] <= 30'b000000010000000000111111000000
                ;mem[3166] <= 30'b000000010000000000111111010000
                ;mem[3167] <= 30'b000000000000000001000011110000
                ;mem[3168] <= 30'b000000000000000001000100000000
                ;mem[3169] <= 30'b000000000000000001000100010000
                ;mem[3170] <= 30'b000000000000000001000100100000
                ;mem[3171] <= 30'b000000000000000001000100110000
                ;mem[3172] <= 30'b000000000000000001000101000000
                ;mem[3173] <= 30'b000000000000000001000101010000
                ;mem[3174] <= 30'b000000000000000001000101100000
                ;mem[3175] <= 30'b000000000000000001001011010000
                ;mem[3176] <= 30'b000000000000000001001011100000
                ;mem[3177] <= 30'b000000000000000001001011110000
                ;mem[3178] <= 30'b000000000000000001001100000000
                ;mem[3179] <= 30'b000000000000000001010010010000
                ;mem[3180] <= 30'b000000000000000001010010100000
                ;mem[3181] <= 30'b000000000000000001010010110000
                ;mem[3182] <= 30'b000000000000000001010011000000
                ;mem[3183] <= 30'b000000000000000001010011010000
                ;mem[3184] <= 30'b000000000000000001011001100000
                ;mem[3185] <= 30'b000000000000000001011001110000
                ;mem[3186] <= 30'b000000000000000001011010000000
                ;mem[3187] <= 30'b000000000000000000100111010000
                ;mem[3188] <= 30'b000000000000000000100111100000
                ;mem[3189] <= 30'b000000000000000000100111110000
                ;mem[3190] <= 30'b000000000000000000101000000000
                ;mem[3191] <= 30'b000000000000000000101000010000
                ;mem[3192] <= 30'b000000000000000000101000100000
                ;mem[3193] <= 30'b000000000000000000101000110000
                ;mem[3194] <= 30'b000000000000000000101101100000
                ;mem[3195] <= 30'b000000000000000000101101110000
                ;mem[3196] <= 30'b000000000000000000101110000000
                ;mem[3197] <= 30'b000000000000000000101110010000
                ;mem[3198] <= 30'b000000000000000000101110100000
                ;mem[3199] <= 30'b000000000000000000101110110000
                ;mem[3200] <= 30'b000000000000000000101111100000
                ;mem[3201] <= 30'b000000000000000000101111110000
                ;mem[3202] <= 30'b000000000000000000110000000000
                ;mem[3203] <= 30'b000000000000000000110011110000
                ;mem[3204] <= 30'b000000000000000000110100000000
                ;mem[3205] <= 30'b000000000000000000110100010000
                ;mem[3206] <= 30'b000000000000000000110100100000
                ;mem[3207] <= 30'b000000000000000000110100110000
                ;mem[3208] <= 30'b000000000000000000110101000000
                ;mem[3209] <= 30'b000000000000000000110110110000
                ;mem[3210] <= 30'b000000000000000000111010110000
                ;mem[3211] <= 30'b000000000000000000111011000000
                ;mem[3212] <= 30'b000000000000000000111011010000
                ;mem[3213] <= 30'b000000001000000000000001100000
                ;mem[3214] <= 30'b000000001000000000000001110000
                ;mem[3215] <= 30'b000000001000000000000010000000
                ;mem[3216] <= 30'b000000001000000000000010010000
                ;mem[3217] <= 30'b000000001000000000000010100000
                ;mem[3218] <= 30'b000000001000000000000010110000
                ;mem[3219] <= 30'b000000001000000000000011100000
                ;mem[3220] <= 30'b000000001000000000000011110000
                ;mem[3221] <= 30'b000000001000000000000100000000
                ;mem[3222] <= 30'b000000001000000000000111110000
                ;mem[3223] <= 30'b000000001000000000001000000000
                ;mem[3224] <= 30'b000000001000000000001000010000
                ;mem[3225] <= 30'b000000001000000000001000100000
                ;mem[3226] <= 30'b000000001000000000001000110000
                ;mem[3227] <= 30'b000000001000000000001001000000
                ;mem[3228] <= 30'b000000001000000000001010110000
                ;mem[3229] <= 30'b000000001000000000001110110000
                ;mem[3230] <= 30'b000000001000000000001111000000
                ;mem[3231] <= 30'b000000001000000000001111010000
                ;mem[3232] <= 30'b000000001000000000010101110000
                ;mem[3233] <= 30'b000000001000000000010110000000
                ;mem[3234] <= 30'b000000001000000000011100110000
                ;mem[3235] <= 30'b000000001000000000011101000000
                ;mem[3236] <= 30'b000000001000000000100011100000
                ;mem[3237] <= 30'b000000001000000000100011110000
                ;mem[3238] <= 30'b000000001000000000100100000000
                ;mem[3239] <= 30'b000000001000000000101010100000
                ;mem[3240] <= 30'b000000001000000000101010110000
                ;mem[3241] <= 30'b000000001000000000110001100000
                ;mem[3242] <= 30'b000000001000000000110001110000
                ;mem[3243] <= 30'b000000001000000000111000100000
                ;mem[3244] <= 30'b000000001000000000111000110000
                ;mem[3245] <= 30'b000000001000000000111111100000
                ;mem[3246] <= 30'b000000001000000000111111110000
                ;mem[3247] <= 30'b000000010000000000000101100000
                ;mem[3248] <= 30'b000000010000000000000101110000
                ;mem[3249] <= 30'b000000010000000000001100100000
                ;mem[3250] <= 30'b000000010000000000001100110000
                ;mem[3251] <= 30'b000000010000000000010011100000
                ;mem[3252] <= 30'b000000010000000000010011110000
                ;mem[3253] <= 30'b000000010000000000010100000000
                ;mem[3254] <= 30'b000000010000000000010100010000
                ;mem[3255] <= 30'b000000010000000000010100100000
                ;mem[3256] <= 30'b000000010000000000010100110000
                ;mem[3257] <= 30'b000000010000000000010101000000
                ;mem[3258] <= 30'b000000010000000000011010100000
                ;mem[3259] <= 30'b000000010000000000011010110000
                ;mem[3260] <= 30'b000000010000000000011011000000
                ;mem[3261] <= 30'b000000010000000000011011010000
                ;mem[3262] <= 30'b000000010000000000011011100000
                ;mem[3263] <= 30'b000000010000000000011011110000
                ;mem[3264] <= 30'b000000010000000000011100000000
                ;mem[3265] <= 30'b000000010000000000011100010000
                ;mem[3266] <= 30'b000000010000000000011100100000
                ;mem[3267] <= 30'b000000010000000000100011010000
                ;mem[3268] <= 30'b000000010000000000100011100000
                ;mem[3269] <= 30'b000000010000000000101010010000
                ;mem[3270] <= 30'b000000010000000000101010100000
                ;mem[3271] <= 30'b000000010000000000110001000000
                ;mem[3272] <= 30'b000000010000000000110001010000
                ;mem[3273] <= 30'b000000010000000000110001100000
                ;mem[3274] <= 30'b000000010000000000110111100000
                ;mem[3275] <= 30'b000000010000000000110111110000
                ;mem[3276] <= 30'b000000010000000000111000000000
                ;mem[3277] <= 30'b000000010000000000111000010000
                ;mem[3278] <= 30'b000000010000000000111110000000
                ;mem[3279] <= 30'b000000010000000000111110010000
                ;mem[3280] <= 30'b000000010000000000111110100000
                ;mem[3281] <= 30'b000000010000000000111110110000
                ;mem[3282] <= 30'b000000000000000001000101000000
                ;mem[3283] <= 30'b000000000000000001000101010000
                ;mem[3284] <= 30'b000000000000000001000101100000
                ;mem[3285] <= 30'b000000000000000001001011100000
                ;mem[3286] <= 30'b000000000000000001001011110000
                ;mem[3287] <= 30'b000000000000000001001100000000
                ;mem[3288] <= 30'b000000000000000001001100010000
                ;mem[3289] <= 30'b000000000000000001010010000000
                ;mem[3290] <= 30'b000000000000000001010010010000
                ;mem[3291] <= 30'b000000000000000001010010100000
                ;mem[3292] <= 30'b000000000000000001010010110000
                ;mem[3293] <= 30'b000000000000000001011000010000
                ;mem[3294] <= 30'b000000000000000001011000100000
                ;mem[3295] <= 30'b000000000000000001011000110000
                ;mem[3296] <= 30'b000000000000000001011001000000
                ;mem[3297] <= 30'b000000000000000001011001010000
                ;mem[3298] <= 30'b000000000000000001011001100000
                ;mem[3299] <= 30'b000000000000000001011110110000
                ;mem[3300] <= 30'b000000000000000001011111000000
                ;mem[3301] <= 30'b000000000000000001011111010000
                ;mem[3302] <= 30'b000000000000000001011111100000
                ;mem[3303] <= 30'b000000000000000001011111110000
                ;mem[3304] <= 30'b000000000000000001100000000000
                ;mem[3305] <= 30'b000000000000000001100110000000
                ;mem[3306] <= 30'b000000000000000001100110010000
                ;mem[3307] <= 30'b000000000000000000100101110000
                ;mem[3308] <= 30'b000000000000000000101100110000
                ;mem[3309] <= 30'b000000000000000000110011100000
                ;mem[3310] <= 30'b000000000000000000110011110000
                ;mem[3311] <= 30'b000000000000000000110101000000
                ;mem[3312] <= 30'b000000000000000000111010100000
                ;mem[3313] <= 30'b000000000000000000111100000000
                ;mem[3314] <= 30'b000000000000000000111100010000
                ;mem[3315] <= 30'b000000001000000000000000110000
                ;mem[3316] <= 30'b000000001000000000000111100000
                ;mem[3317] <= 30'b000000001000000000000111110000
                ;mem[3318] <= 30'b000000001000000000001001000000
                ;mem[3319] <= 30'b000000001000000000001110100000
                ;mem[3320] <= 30'b000000001000000000010000000000
                ;mem[3321] <= 30'b000000001000000000010000010000
                ;mem[3322] <= 30'b000000001000000000010101010000
                ;mem[3323] <= 30'b000000001000000000010111010000
                ;mem[3324] <= 30'b000000001000000000011100010000
                ;mem[3325] <= 30'b000000001000000000011110010000
                ;mem[3326] <= 30'b000000001000000000100011010000
                ;mem[3327] <= 30'b000000001000000000100101000000
                ;mem[3328] <= 30'b000000001000000000100101010000
                ;mem[3329] <= 30'b000000001000000000101010000000
                ;mem[3330] <= 30'b000000001000000000101100000000
                ;mem[3331] <= 30'b000000001000000000101100010000
                ;mem[3332] <= 30'b000000001000000000110001000000
                ;mem[3333] <= 30'b000000001000000000110011000000
                ;mem[3334] <= 30'b000000001000000000110011010000
                ;mem[3335] <= 30'b000000001000000000110111110000
                ;mem[3336] <= 30'b000000001000000000111000000000
                ;mem[3337] <= 30'b000000001000000000111010000000
                ;mem[3338] <= 30'b000000001000000000111010010000
                ;mem[3339] <= 30'b000000001000000000111110110000
                ;mem[3340] <= 30'b000000001000000000111111000000
                ;mem[3341] <= 30'b000000001000000000111111010000
                ;mem[3342] <= 30'b000000010000000000000000000000
                ;mem[3343] <= 30'b000000010000000000000000010000
                ;mem[3344] <= 30'b000000010000000000000101000000
                ;mem[3345] <= 30'b000000010000000000000111000000
                ;mem[3346] <= 30'b000000010000000000000111010000
                ;mem[3347] <= 30'b000000010000000000001011110000
                ;mem[3348] <= 30'b000000010000000000001100000000
                ;mem[3349] <= 30'b000000010000000000001110000000
                ;mem[3350] <= 30'b000000010000000000001110010000
                ;mem[3351] <= 30'b000000010000000000010010110000
                ;mem[3352] <= 30'b000000010000000000010011000000
                ;mem[3353] <= 30'b000000010000000000010011010000
                ;mem[3354] <= 30'b000000010000000000010101010000
                ;mem[3355] <= 30'b000000010000000000011010010000
                ;mem[3356] <= 30'b000000010000000000011010100000
                ;mem[3357] <= 30'b000000010000000000011010110000
                ;mem[3358] <= 30'b000000010000000000011011000000
                ;mem[3359] <= 30'b000000010000000000011011010000
                ;mem[3360] <= 30'b000000010000000000011011100000
                ;mem[3361] <= 30'b000000010000000000011011110000
                ;mem[3362] <= 30'b000000010000000000011100000000
                ;mem[3363] <= 30'b000000010000000000011100010000
                ;mem[3364] <= 30'b000000010000000000011100100000
                ;mem[3365] <= 30'b000000010000000000011100110000
                ;mem[3366] <= 30'b000000010000000000100011000000
                ;mem[3367] <= 30'b000000010000000000100011010000
                ;mem[3368] <= 30'b000000010000000000101010000000
                ;mem[3369] <= 30'b000000010000000000101010010000
                ;mem[3370] <= 30'b000000010000000000110001000000
                ;mem[3371] <= 30'b000000010000000000110001010000
                ;mem[3372] <= 30'b000000010000000000111000010000
                ;mem[3373] <= 30'b000000010000000000111111010000
                ;mem[3374] <= 30'b000000000000000001000101000000
                ;mem[3375] <= 30'b000000000000000001000101010000
                ;mem[3376] <= 30'b000000000000000001001100010000
                ;mem[3377] <= 30'b000000000000000001010011010000
                ;mem[3378] <= 30'b000000000000000001011010010000
                ;mem[3379] <= 30'b000000000000000001100001010000
                ;mem[3380] <= 30'b000000000000000001100001100000
                ;mem[3381] <= 30'b000000000000000001101000100000
                ;mem[3382] <= 30'b000000000000000000011111110000
                ;mem[3383] <= 30'b000000000000000000100110100000
                ;mem[3384] <= 30'b000000000000000000100110110000
                ;mem[3385] <= 30'b000000000000000000100111000000
                ;mem[3386] <= 30'b000000000000000000100111010000
                ;mem[3387] <= 30'b000000000000000000100111100000
                ;mem[3388] <= 30'b000000000000000000100111110000
                ;mem[3389] <= 30'b000000000000000000101000000000
                ;mem[3390] <= 30'b000000000000000000101101100000
                ;mem[3391] <= 30'b000000000000000000101101110000
                ;mem[3392] <= 30'b000000000000000000101110000000
                ;mem[3393] <= 30'b000000000000000000101110010000
                ;mem[3394] <= 30'b000000000000000000101110100000
                ;mem[3395] <= 30'b000000000000000000101110110000
                ;mem[3396] <= 30'b000000000000000000101111000000
                ;mem[3397] <= 30'b000000000000000000101111010000
                ;mem[3398] <= 30'b000000000000000000110011010000
                ;mem[3399] <= 30'b000000000000000000110011100000
                ;mem[3400] <= 30'b000000000000000000110011110000
                ;mem[3401] <= 30'b000000000000000000110100100000
                ;mem[3402] <= 30'b000000000000000000110100110000
                ;mem[3403] <= 30'b000000000000000000110101000000
                ;mem[3404] <= 30'b000000000000000000110101010000
                ;mem[3405] <= 30'b000000000000000000110101100000
                ;mem[3406] <= 30'b000000000000000000110101110000
                ;mem[3407] <= 30'b000000000000000000110110000000
                ;mem[3408] <= 30'b000000000000000000110110010000
                ;mem[3409] <= 30'b000000000000000000111010000000
                ;mem[3410] <= 30'b000000000000000000111010010000
                ;mem[3411] <= 30'b000000000000000000111010100000
                ;mem[3412] <= 30'b000000000000000000111010110000
                ;mem[3413] <= 30'b000000000000000000111011000000
                ;mem[3414] <= 30'b000000000000000000111011110000
                ;mem[3415] <= 30'b000000000000000000111100000000
                ;mem[3416] <= 30'b000000000000000000111100010000
                ;mem[3417] <= 30'b000000000000000000111100100000
                ;mem[3418] <= 30'b000000000000000000111100110000
                ;mem[3419] <= 30'b000000000000000000111101000000
                ;mem[3420] <= 30'b000000000000000000111101010000
                ;mem[3421] <= 30'b000000000000000000111101100000
                ;mem[3422] <= 30'b000000001000000000000001100000
                ;mem[3423] <= 30'b000000001000000000000001110000
                ;mem[3424] <= 30'b000000001000000000000010000000
                ;mem[3425] <= 30'b000000001000000000000010010000
                ;mem[3426] <= 30'b000000001000000000000010100000
                ;mem[3427] <= 30'b000000001000000000000010110000
                ;mem[3428] <= 30'b000000001000000000000011000000
                ;mem[3429] <= 30'b000000001000000000000011010000
                ;mem[3430] <= 30'b000000001000000000000111010000
                ;mem[3431] <= 30'b000000001000000000000111100000
                ;mem[3432] <= 30'b000000001000000000000111110000
                ;mem[3433] <= 30'b000000001000000000001000100000
                ;mem[3434] <= 30'b000000001000000000001000110000
                ;mem[3435] <= 30'b000000001000000000001001000000
                ;mem[3436] <= 30'b000000001000000000001001010000
                ;mem[3437] <= 30'b000000001000000000001001100000
                ;mem[3438] <= 30'b000000001000000000001001110000
                ;mem[3439] <= 30'b000000001000000000001010000000
                ;mem[3440] <= 30'b000000001000000000001010010000
                ;mem[3441] <= 30'b000000001000000000001110000000
                ;mem[3442] <= 30'b000000001000000000001110010000
                ;mem[3443] <= 30'b000000001000000000001110100000
                ;mem[3444] <= 30'b000000001000000000001110110000
                ;mem[3445] <= 30'b000000001000000000001111000000
                ;mem[3446] <= 30'b000000001000000000001111110000
                ;mem[3447] <= 30'b000000001000000000010000000000
                ;mem[3448] <= 30'b000000001000000000010000010000
                ;mem[3449] <= 30'b000000001000000000010000100000
                ;mem[3450] <= 30'b000000001000000000010000110000
                ;mem[3451] <= 30'b000000001000000000010001000000
                ;mem[3452] <= 30'b000000001000000000010001010000
                ;mem[3453] <= 30'b000000001000000000010001100000
                ;mem[3454] <= 30'b000000001000000000010100110000
                ;mem[3455] <= 30'b000000001000000000010101000000
                ;mem[3456] <= 30'b000000001000000000010101010000
                ;mem[3457] <= 30'b000000001000000000010101100000
                ;mem[3458] <= 30'b000000001000000000010101110000
                ;mem[3459] <= 30'b000000001000000000010110000000
                ;mem[3460] <= 30'b000000001000000000010111000000
                ;mem[3461] <= 30'b000000001000000000010111010000
                ;mem[3462] <= 30'b000000001000000000010111100000
                ;mem[3463] <= 30'b000000001000000000010111110000
                ;mem[3464] <= 30'b000000001000000000011000000000
                ;mem[3465] <= 30'b000000001000000000011000010000
                ;mem[3466] <= 30'b000000001000000000011000100000
                ;mem[3467] <= 30'b000000001000000000011011100000
                ;mem[3468] <= 30'b000000001000000000011011110000
                ;mem[3469] <= 30'b000000001000000000011100000000
                ;mem[3470] <= 30'b000000001000000000011100010000
                ;mem[3471] <= 30'b000000001000000000011100100000
                ;mem[3472] <= 30'b000000001000000000011100110000
                ;mem[3473] <= 30'b000000001000000000011101000000
                ;mem[3474] <= 30'b000000001000000000011111000000
                ;mem[3475] <= 30'b000000001000000000011111010000
                ;mem[3476] <= 30'b000000001000000000011111100000
                ;mem[3477] <= 30'b000000001000000000011111110000
                ;mem[3478] <= 30'b000000001000000000100010100000
                ;mem[3479] <= 30'b000000001000000000100010110000
                ;mem[3480] <= 30'b000000001000000000100011000000
                ;mem[3481] <= 30'b000000001000000000100011010000
                ;mem[3482] <= 30'b000000001000000000100011100000
                ;mem[3483] <= 30'b000000001000000000100011110000
                ;mem[3484] <= 30'b000000001000000000100100000000
                ;mem[3485] <= 30'b000000001000000000100110010000
                ;mem[3486] <= 30'b000000001000000000100110100000
                ;mem[3487] <= 30'b000000001000000000100110110000
                ;mem[3488] <= 30'b000000001000000000101001100000
                ;mem[3489] <= 30'b000000001000000000101001110000
                ;mem[3490] <= 30'b000000001000000000101010000000
                ;mem[3491] <= 30'b000000001000000000101010010000
                ;mem[3492] <= 30'b000000001000000000101010100000
                ;mem[3493] <= 30'b000000001000000000101010110000
                ;mem[3494] <= 30'b000000001000000000101101010000
                ;mem[3495] <= 30'b000000001000000000101101100000
                ;mem[3496] <= 30'b000000001000000000101101110000
                ;mem[3497] <= 30'b000000001000000000110000010000
                ;mem[3498] <= 30'b000000001000000000110000100000
                ;mem[3499] <= 30'b000000001000000000110000110000
                ;mem[3500] <= 30'b000000001000000000110001000000
                ;mem[3501] <= 30'b000000001000000000110001010000
                ;mem[3502] <= 30'b000000001000000000110001100000
                ;mem[3503] <= 30'b000000001000000000110001110000
                ;mem[3504] <= 30'b000000001000000000110100000000
                ;mem[3505] <= 30'b000000001000000000110100010000
                ;mem[3506] <= 30'b000000001000000000110100100000
                ;mem[3507] <= 30'b000000001000000000110100110000
                ;mem[3508] <= 30'b000000001000000000110111010000
                ;mem[3509] <= 30'b000000001000000000110111100000
                ;mem[3510] <= 30'b000000001000000000110111110000
                ;mem[3511] <= 30'b000000001000000000111000000000
                ;mem[3512] <= 30'b000000001000000000111000010000
                ;mem[3513] <= 30'b000000001000000000111000100000
                ;mem[3514] <= 30'b000000001000000000111011000000
                ;mem[3515] <= 30'b000000001000000000111011010000
                ;mem[3516] <= 30'b000000001000000000111011100000
                ;mem[3517] <= 30'b000000001000000000111011110000
                ;mem[3518] <= 30'b000000001000000000111110010000
                ;mem[3519] <= 30'b000000001000000000111110100000
                ;mem[3520] <= 30'b000000001000000000111110110000
                ;mem[3521] <= 30'b000000001000000000111111000000
                ;mem[3522] <= 30'b000000001000000000111111010000
                ;mem[3523] <= 30'b000000010000000000000001010000
                ;mem[3524] <= 30'b000000010000000000000001100000
                ;mem[3525] <= 30'b000000010000000000000001110000
                ;mem[3526] <= 30'b000000010000000000000100010000
                ;mem[3527] <= 30'b000000010000000000000100100000
                ;mem[3528] <= 30'b000000010000000000000100110000
                ;mem[3529] <= 30'b000000010000000000000101000000
                ;mem[3530] <= 30'b000000010000000000000101010000
                ;mem[3531] <= 30'b000000010000000000000101100000
                ;mem[3532] <= 30'b000000010000000000000101110000
                ;mem[3533] <= 30'b000000010000000000001000000000
                ;mem[3534] <= 30'b000000010000000000001000010000
                ;mem[3535] <= 30'b000000010000000000001000100000
                ;mem[3536] <= 30'b000000010000000000001000110000
                ;mem[3537] <= 30'b000000010000000000001011010000
                ;mem[3538] <= 30'b000000010000000000001011100000
                ;mem[3539] <= 30'b000000010000000000001011110000
                ;mem[3540] <= 30'b000000010000000000001100000000
                ;mem[3541] <= 30'b000000010000000000001100010000
                ;mem[3542] <= 30'b000000010000000000001100100000
                ;mem[3543] <= 30'b000000010000000000001111000000
                ;mem[3544] <= 30'b000000010000000000001111010000
                ;mem[3545] <= 30'b000000010000000000001111100000
                ;mem[3546] <= 30'b000000010000000000001111110000
                ;mem[3547] <= 30'b000000010000000000010010010000
                ;mem[3548] <= 30'b000000010000000000010010100000
                ;mem[3549] <= 30'b000000010000000000010010110000
                ;mem[3550] <= 30'b000000010000000000010011000000
                ;mem[3551] <= 30'b000000010000000000010011010000
                ;mem[3552] <= 30'b000000010000000000010101100000
                ;mem[3553] <= 30'b000000010000000000010101110000
                ;mem[3554] <= 30'b000000010000000000010110000000
                ;mem[3555] <= 30'b000000010000000000010110010000
                ;mem[3556] <= 30'b000000010000000000010110100000
                ;mem[3557] <= 30'b000000010000000000010110110000
                ;mem[3558] <= 30'b000000010000000000011001010000
                ;mem[3559] <= 30'b000000010000000000011001100000
                ;mem[3560] <= 30'b000000010000000000011001110000
                ;mem[3561] <= 30'b000000010000000000011010000000
                ;mem[3562] <= 30'b000000010000000000011010010000
                ;mem[3563] <= 30'b000000010000000000011100000000
                ;mem[3564] <= 30'b000000010000000000011100010000
                ;mem[3565] <= 30'b000000010000000000011100100000
                ;mem[3566] <= 30'b000000010000000000011100110000
                ;mem[3567] <= 30'b000000010000000000011101000000
                ;mem[3568] <= 30'b000000010000000000011101010000
                ;mem[3569] <= 30'b000000010000000000011101100000
                ;mem[3570] <= 30'b000000010000000000100000010000
                ;mem[3571] <= 30'b000000010000000000100000100000
                ;mem[3572] <= 30'b000000010000000000100000110000
                ;mem[3573] <= 30'b000000010000000000100001000000
                ;mem[3574] <= 30'b000000010000000000100001010000
                ;mem[3575] <= 30'b000000010000000000100010010000
                ;mem[3576] <= 30'b000000010000000000100010100000
                ;mem[3577] <= 30'b000000010000000000100010110000
                ;mem[3578] <= 30'b000000010000000000100011000000
                ;mem[3579] <= 30'b000000010000000000100011010000
                ;mem[3580] <= 30'b000000010000000000100011100000
                ;mem[3581] <= 30'b000000010000000000100011110000
                ;mem[3582] <= 30'b000000010000000000100100000000
                ;mem[3583] <= 30'b000000010000000000100100010000
                ;mem[3584] <= 30'b000000010000000000100111010000
                ;mem[3585] <= 30'b000000010000000000100111100000
                ;mem[3586] <= 30'b000000010000000000100111110000
                ;mem[3587] <= 30'b000000010000000000101000000000
                ;mem[3588] <= 30'b000000010000000000101000010000
                ;mem[3589] <= 30'b000000010000000000101000100000
                ;mem[3590] <= 30'b000000010000000000101000110000
                ;mem[3591] <= 30'b000000010000000000101001000000
                ;mem[3592] <= 30'b000000010000000000101001010000
                ;mem[3593] <= 30'b000000010000000000101001100000
                ;mem[3594] <= 30'b000000010000000000101001110000
                ;mem[3595] <= 30'b000000010000000000101010000000
                ;mem[3596] <= 30'b000000010000000000101010010000
                ;mem[3597] <= 30'b000000010000000000101010100000
                ;mem[3598] <= 30'b000000010000000000101010110000
                ;mem[3599] <= 30'b000000010000000000101011000000
                ;mem[3600] <= 30'b000000010000000000101011010000
                ;mem[3601] <= 30'b000000010000000000101110100000
                ;mem[3602] <= 30'b000000010000000000101110110000
                ;mem[3603] <= 30'b000000010000000000101111000000
                ;mem[3604] <= 30'b000000010000000000101111010000
                ;mem[3605] <= 30'b000000010000000000101111100000
                ;mem[3606] <= 30'b000000010000000000101111110000
                ;mem[3607] <= 30'b000000010000000000110000000000
                ;mem[3608] <= 30'b000000010000000000110000010000
                ;mem[3609] <= 30'b000000010000000000110000100000
                ;mem[3610] <= 30'b000000010000000000110000110000
                ;mem[3611] <= 30'b000000010000000000110001000000
                ;mem[3612] <= 30'b000000010000000000110001010000
                ;mem[3613] <= 30'b000000010000000000110001100000
                ;mem[3614] <= 30'b000000010000000000110001110000
                ;mem[3615] <= 30'b000000010000000000110010000000
                ;mem[3616] <= 30'b000000010000000000110101100000
                ;mem[3617] <= 30'b000000010000000000110101110000
                ;mem[3618] <= 30'b000000010000000000110110000000
                ;mem[3619] <= 30'b000000010000000000110110010000
                ;mem[3620] <= 30'b000000010000000000110110100000
                ;mem[3621] <= 30'b000000010000000000110110110000
                ;mem[3622] <= 30'b000000010000000000110111000000
                ;mem[3623] <= 30'b000000010000000000110111010000
                ;mem[3624] <= 30'b000000010000000000110111100000
                ;mem[3625] <= 30'b000000010000000000110111110000
                ;mem[3626] <= 30'b000000010000000000111000000000
                ;mem[3627] <= 30'b000000010000000000111000010000
                ;mem[3628] <= 30'b000000010000000000111000100000
                ;mem[3629] <= 30'b000000010000000000111100110000
                ;mem[3630] <= 30'b000000010000000000111101000000
                ;mem[3631] <= 30'b000000010000000000111101010000
                ;mem[3632] <= 30'b000000010000000000111101100000
                ;mem[3633] <= 30'b000000010000000000111101110000
                ;mem[3634] <= 30'b000000010000000000111110000000
                ;mem[3635] <= 30'b000000010000000000111110010000
                ;mem[3636] <= 30'b000000010000000000111110100000
                ;mem[3637] <= 30'b000000010000000000111110110000
                ;mem[3638] <= 30'b000000010000000000111111000000
                ;mem[3639] <= 30'b000000010000000000111111010000
                ;mem[3640] <= 30'b000000000000000001000010100000
                ;mem[3641] <= 30'b000000000000000001000010110000
                ;mem[3642] <= 30'b000000000000000001000011000000
                ;mem[3643] <= 30'b000000000000000001000011010000
                ;mem[3644] <= 30'b000000000000000001000011100000
                ;mem[3645] <= 30'b000000000000000001000011110000
                ;mem[3646] <= 30'b000000000000000001000100000000
                ;mem[3647] <= 30'b000000000000000001000100010000
                ;mem[3648] <= 30'b000000000000000001000100100000
                ;mem[3649] <= 30'b000000000000000001000100110000
                ;mem[3650] <= 30'b000000000000000001000101000000
                ;mem[3651] <= 30'b000000000000000001000101010000
                ;mem[3652] <= 30'b000000000000000001000101100000
                ;mem[3653] <= 30'b000000000000000001000101110000
                ;mem[3654] <= 30'b000000000000000001000110000000
                ;mem[3655] <= 30'b000000000000000001001001100000
                ;mem[3656] <= 30'b000000000000000001001001110000
                ;mem[3657] <= 30'b000000000000000001001010000000
                ;mem[3658] <= 30'b000000000000000001001010010000
                ;mem[3659] <= 30'b000000000000000001001010100000
                ;mem[3660] <= 30'b000000000000000001001010110000
                ;mem[3661] <= 30'b000000000000000001001011000000
                ;mem[3662] <= 30'b000000000000000001001011010000
                ;mem[3663] <= 30'b000000000000000001001011100000
                ;mem[3664] <= 30'b000000000000000001001011110000
                ;mem[3665] <= 30'b000000000000000001001100000000
                ;mem[3666] <= 30'b000000000000000001001100010000
                ;mem[3667] <= 30'b000000000000000001001100100000
                ;mem[3668] <= 30'b000000000000000001010000110000
                ;mem[3669] <= 30'b000000000000000001010001000000
                ;mem[3670] <= 30'b000000000000000001010001010000
                ;mem[3671] <= 30'b000000000000000001010001100000
                ;mem[3672] <= 30'b000000000000000001010001110000
                ;mem[3673] <= 30'b000000000000000001010010000000
                ;mem[3674] <= 30'b000000000000000001010010010000
                ;mem[3675] <= 30'b000000000000000001010010100000
                ;mem[3676] <= 30'b000000000000000001010010110000
                ;mem[3677] <= 30'b000000000000000001010011000000
                ;mem[3678] <= 30'b000000000000000001010011010000
                ;mem[3679] <= 30'b000000000000000001011000000000
                ;mem[3680] <= 30'b000000000000000001011000010000
                ;mem[3681] <= 30'b000000000000000001011000100000
                ;mem[3682] <= 30'b000000000000000001011000110000
                ;mem[3683] <= 30'b000000000000000001011001000000
                ;mem[3684] <= 30'b000000000000000001011001010000
                ;mem[3685] <= 30'b000000000000000001011001100000
                ;mem[3686] <= 30'b000000000000000001011001110000
                ;mem[3687] <= 30'b000000000000000001011111100000
                ;mem[3688] <= 30'b000000000000000001011111110000
                ;mem[3689] <= 30'b000000000000000001100000000000
                ;mem[3690] <= 30'b000000000000000000111011000000
                ;mem[3691] <= 30'b000000000000000000111011010000
                ;mem[3692] <= 30'b000000000000000000111011100000
                ;mem[3693] <= 30'b000000000000000000111011110000
                ;mem[3694] <= 30'b000000000000000000111100000000
                ;mem[3695] <= 30'b000000000000000000111100010000
                ;mem[3696] <= 30'b000000001000000000001111000000
                ;mem[3697] <= 30'b000000001000000000001111010000
                ;mem[3698] <= 30'b000000001000000000001111100000
                ;mem[3699] <= 30'b000000001000000000001111110000
                ;mem[3700] <= 30'b000000001000000000010000000000
                ;mem[3701] <= 30'b000000001000000000010000010000
                ;mem[3702] <= 30'b000000001000000000010100100000
                ;mem[3703] <= 30'b000000001000000000010101100000
                ;mem[3704] <= 30'b000000001000000000010101110000
                ;mem[3705] <= 30'b000000001000000000010110000000
                ;mem[3706] <= 30'b000000001000000000010110010000
                ;mem[3707] <= 30'b000000001000000000010110100000
                ;mem[3708] <= 30'b000000001000000000010110110000
                ;mem[3709] <= 30'b000000001000000000010111000000
                ;mem[3710] <= 30'b000000001000000000010111010000
                ;mem[3711] <= 30'b000000001000000000010111100000
                ;mem[3712] <= 30'b000000001000000000011011010000
                ;mem[3713] <= 30'b000000001000000000011011100000
                ;mem[3714] <= 30'b000000001000000000011011110000
                ;mem[3715] <= 30'b000000001000000000011100000000
                ;mem[3716] <= 30'b000000001000000000011100010000
                ;mem[3717] <= 30'b000000001000000000011100100000
                ;mem[3718] <= 30'b000000001000000000011110000000
                ;mem[3719] <= 30'b000000001000000000011110010000
                ;mem[3720] <= 30'b000000001000000000011110100000
                ;mem[3721] <= 30'b000000001000000000100010010000
                ;mem[3722] <= 30'b000000001000000000100010100000
                ;mem[3723] <= 30'b000000001000000000100010110000
                ;mem[3724] <= 30'b000000001000000000100011000000
                ;mem[3725] <= 30'b000000001000000000100101010000
                ;mem[3726] <= 30'b000000001000000000100101100000
                ;mem[3727] <= 30'b000000001000000000100101110000
                ;mem[3728] <= 30'b000000001000000000101001010000
                ;mem[3729] <= 30'b000000001000000000101100010000
                ;mem[3730] <= 30'b000000001000000000101100100000
                ;mem[3731] <= 30'b000000001000000000101100110000
                ;mem[3732] <= 30'b000000001000000000110011010000
                ;mem[3733] <= 30'b000000001000000000110011100000
                ;mem[3734] <= 30'b000000001000000000110011110000
                ;mem[3735] <= 30'b000000001000000000111010100000
                ;mem[3736] <= 30'b000000001000000000111010110000
                ;mem[3737] <= 30'b000000010000000000000000010000
                ;mem[3738] <= 30'b000000010000000000000000100000
                ;mem[3739] <= 30'b000000010000000000000000110000
                ;mem[3740] <= 30'b000000010000000000000111010000
                ;mem[3741] <= 30'b000000010000000000000111100000
                ;mem[3742] <= 30'b000000010000000000000111110000
                ;mem[3743] <= 30'b000000010000000000001110100000
                ;mem[3744] <= 30'b000000010000000000001110110000
                ;mem[3745] <= 30'b000000010000000000010101100000
                ;mem[3746] <= 30'b000000010000000000010101110000
                ;mem[3747] <= 30'b000000010000000000011100010000
                ;mem[3748] <= 30'b000000010000000000011100100000
                ;mem[3749] <= 30'b000000010000000000100011010000
                ;mem[3750] <= 30'b000000010000000000100011100000
                ;mem[3751] <= 30'b000000010000000000101010010000
                ;mem[3752] <= 30'b000000010000000000101010100000
                ;mem[3753] <= 30'b000000010000000000110001010000
                ;mem[3754] <= 30'b000000010000000000111000010000
                ;mem[3755] <= 30'b000000010000000000111111000000
                ;mem[3756] <= 30'b000000010000000000111111010000
                ;mem[3757] <= 30'b000000000000000001000101010000
                ;mem[3758] <= 30'b000000000000000001001100010000
                ;mem[3759] <= 30'b000000000000000001010011000000
                ;mem[3760] <= 30'b000000000000000001010011010000
                ;mem[3761] <= 30'b000000000000000001011010000000
                ;mem[3762] <= 30'b000000000000000001011010010000
                ;mem[3763] <= 30'b000000000000000001100001000000
                ;mem[3764] <= 30'b000000000000000001100001010000
                ;mem[3765] <= 30'b000000000000000001101000000000
                ;mem[3766] <= 30'b000000000000000001101110110000
                ;mem[3767] <= 30'b000000000000000001101111000000
                ;mem[3768] <= 30'b000000000000000001110101110000
                ;mem[3769] <= 30'b000000000000000001110110000000
                ;mem[3770] <= 30'b000000000000000001111100110000
                ;mem[3771] <= 30'b000000000000000000100110000000
                ;mem[3772] <= 30'b000000000000000000101101000000
                ;mem[3773] <= 30'b000000000000000000101101010000
                ;mem[3774] <= 30'b000000000000000000101110110000
                ;mem[3775] <= 30'b000000000000000000101111000000
                ;mem[3776] <= 30'b000000000000000000110011110000
                ;mem[3777] <= 30'b000000000000000000110100000000
                ;mem[3778] <= 30'b000000000000000000110101110000
                ;mem[3779] <= 30'b000000000000000000110110000000
                ;mem[3780] <= 30'b000000000000000000111010110000
                ;mem[3781] <= 30'b000000000000000000111011000000
                ;mem[3782] <= 30'b000000000000000000111100110000
                ;mem[3783] <= 30'b000000000000000000111101000000
                ;mem[3784] <= 30'b000000001000000000000001000000
                ;mem[3785] <= 30'b000000001000000000000001010000
                ;mem[3786] <= 30'b000000001000000000000010110000
                ;mem[3787] <= 30'b000000001000000000000011000000
                ;mem[3788] <= 30'b000000001000000000000111110000
                ;mem[3789] <= 30'b000000001000000000001000000000
                ;mem[3790] <= 30'b000000001000000000001001110000
                ;mem[3791] <= 30'b000000001000000000001010000000
                ;mem[3792] <= 30'b000000001000000000001110110000
                ;mem[3793] <= 30'b000000001000000000001111000000
                ;mem[3794] <= 30'b000000001000000000010000110000
                ;mem[3795] <= 30'b000000001000000000010001000000
                ;mem[3796] <= 30'b000000001000000000010101100000
                ;mem[3797] <= 30'b000000001000000000010101110000
                ;mem[3798] <= 30'b000000001000000000010110000000
                ;mem[3799] <= 30'b000000001000000000010111100000
                ;mem[3800] <= 30'b000000001000000000010111110000
                ;mem[3801] <= 30'b000000001000000000011100100000
                ;mem[3802] <= 30'b000000001000000000011100110000
                ;mem[3803] <= 30'b000000001000000000011110100000
                ;mem[3804] <= 30'b000000001000000000011110110000
                ;mem[3805] <= 30'b000000001000000000100011010000
                ;mem[3806] <= 30'b000000001000000000100011100000
                ;mem[3807] <= 30'b000000001000000000100101100000
                ;mem[3808] <= 30'b000000001000000000100101110000
                ;mem[3809] <= 30'b000000001000000000101010000000
                ;mem[3810] <= 30'b000000001000000000101010010000
                ;mem[3811] <= 30'b000000001000000000101010100000
                ;mem[3812] <= 30'b000000001000000000101100100000
                ;mem[3813] <= 30'b000000001000000000101100110000
                ;mem[3814] <= 30'b000000001000000000110000110000
                ;mem[3815] <= 30'b000000001000000000110001000000
                ;mem[3816] <= 30'b000000001000000000110001010000
                ;mem[3817] <= 30'b000000001000000000110011100000
                ;mem[3818] <= 30'b000000001000000000110011110000
                ;mem[3819] <= 30'b000000001000000000110111110000
                ;mem[3820] <= 30'b000000001000000000111000000000
                ;mem[3821] <= 30'b000000001000000000111000010000
                ;mem[3822] <= 30'b000000001000000000111000100000
                ;mem[3823] <= 30'b000000001000000000111000110000
                ;mem[3824] <= 30'b000000001000000000111010010000
                ;mem[3825] <= 30'b000000001000000000111010100000
                ;mem[3826] <= 30'b000000001000000000111010110000
                ;mem[3827] <= 30'b000000001000000000111110110000
                ;mem[3828] <= 30'b000000001000000000111111000000
                ;mem[3829] <= 30'b000000001000000000111111010000
                ;mem[3830] <= 30'b000000001000000000111111100000
                ;mem[3831] <= 30'b000000001000000000111111110000
                ;mem[3832] <= 30'b000000010000000000000000100000
                ;mem[3833] <= 30'b000000010000000000000000110000
                ;mem[3834] <= 30'b000000010000000000000100110000
                ;mem[3835] <= 30'b000000010000000000000101000000
                ;mem[3836] <= 30'b000000010000000000000101010000
                ;mem[3837] <= 30'b000000010000000000000111100000
                ;mem[3838] <= 30'b000000010000000000000111110000
                ;mem[3839] <= 30'b000000010000000000001011110000
                ;mem[3840] <= 30'b000000010000000000001100000000
                ;mem[3841] <= 30'b000000010000000000001100010000
                ;mem[3842] <= 30'b000000010000000000001100100000
                ;mem[3843] <= 30'b000000010000000000001100110000
                ;mem[3844] <= 30'b000000010000000000001110010000
                ;mem[3845] <= 30'b000000010000000000001110100000
                ;mem[3846] <= 30'b000000010000000000001110110000
                ;mem[3847] <= 30'b000000010000000000010010110000
                ;mem[3848] <= 30'b000000010000000000010011000000
                ;mem[3849] <= 30'b000000010000000000010011010000
                ;mem[3850] <= 30'b000000010000000000010011100000
                ;mem[3851] <= 30'b000000010000000000010011110000
                ;mem[3852] <= 30'b000000010000000000010100000000
                ;mem[3853] <= 30'b000000010000000000010100010000
                ;mem[3854] <= 30'b000000010000000000010100100000
                ;mem[3855] <= 30'b000000010000000000010100110000
                ;mem[3856] <= 30'b000000010000000000010101000000
                ;mem[3857] <= 30'b000000010000000000010101010000
                ;mem[3858] <= 30'b000000010000000000010101100000
                ;mem[3859] <= 30'b000000010000000000010101110000
                ;mem[3860] <= 30'b000000010000000000011010000000
                ;mem[3861] <= 30'b000000010000000000011010010000
                ;mem[3862] <= 30'b000000010000000000011010100000
                ;mem[3863] <= 30'b000000010000000000011010110000
                ;mem[3864] <= 30'b000000010000000000011011000000
                ;mem[3865] <= 30'b000000010000000000011011010000
                ;mem[3866] <= 30'b000000010000000000011011100000
                ;mem[3867] <= 30'b000000010000000000011011110000
                ;mem[3868] <= 30'b000000010000000000011100000000
                ;mem[3869] <= 30'b000000010000000000011100010000
                ;mem[3870] <= 30'b000000010000000000011100100000
                ;mem[3871] <= 30'b000000010000000000100010010000
                ;mem[3872] <= 30'b000000010000000000100010100000
                ;mem[3873] <= 30'b000000010000000000100011000000
                ;mem[3874] <= 30'b000000010000000000100011010000
                ;mem[3875] <= 30'b000000010000000000100011100000
                ;mem[3876] <= 30'b000000010000000000101010000000
                ;mem[3877] <= 30'b000000010000000000101010010000
                ;mem[3878] <= 30'b000000010000000000101010100000
                ;mem[3879] <= 30'b000000010000000000110001000000
                ;mem[3880] <= 30'b000000010000000000110001010000
                ;mem[3881] <= 30'b000000010000000000110001100000
                ;mem[3882] <= 30'b000000010000000000111000000000
                ;mem[3883] <= 30'b000000010000000000111000010000
                ;mem[3884] <= 30'b000000010000000000111000100000
                ;mem[3885] <= 30'b000000010000000000111111000000
                ;mem[3886] <= 30'b000000010000000000111111010000
                ;mem[3887] <= 30'b000000000000000001000101000000
                ;mem[3888] <= 30'b000000000000000001000101010000
                ;mem[3889] <= 30'b000000000000000001000101100000
                ;mem[3890] <= 30'b000000000000000001001100000000
                ;mem[3891] <= 30'b000000000000000001001100010000
                ;mem[3892] <= 30'b000000000000000001001100100000
                ;mem[3893] <= 30'b000000000000000001010011000000
                ;mem[3894] <= 30'b000000000000000001010011010000
                ;mem[3895] <= 30'b000000000000000001011010000000
                ;mem[3896] <= 30'b000000000000000001011010010000
                ;mem[3897] <= 30'b000000000000000001100001000000
                ;mem[3898] <= 30'b000000000000000001100001010000
                ;mem[3899] <= 30'b000000000000000001101000000000
                ;mem[3900] <= 30'b000000000000000000100101100000
                ;mem[3901] <= 30'b000000000000000000100101110000
                ;mem[3902] <= 30'b000000000000000000100110000000
                ;mem[3903] <= 30'b000000000000000000100110010000
                ;mem[3904] <= 30'b000000000000000000100110100000
                ;mem[3905] <= 30'b000000000000000000100110110000
                ;mem[3906] <= 30'b000000000000000000100111000000
                ;mem[3907] <= 30'b000000000000000000100111010000
                ;mem[3908] <= 30'b000000000000000000101100100000
                ;mem[3909] <= 30'b000000000000000000101100110000
                ;mem[3910] <= 30'b000000000000000000101101000000
                ;mem[3911] <= 30'b000000000000000000101101010000
                ;mem[3912] <= 30'b000000000000000000101101100000
                ;mem[3913] <= 30'b000000000000000000101101110000
                ;mem[3914] <= 30'b000000000000000000101110000000
                ;mem[3915] <= 30'b000000000000000000101110010000
                ;mem[3916] <= 30'b000000000000000000101110100000
                ;mem[3917] <= 30'b000000000000000000110011100000
                ;mem[3918] <= 30'b000000000000000000110011110000
                ;mem[3919] <= 30'b000000000000000000110100000000
                ;mem[3920] <= 30'b000000000000000000110100010000
                ;mem[3921] <= 30'b000000000000000000110100100000
                ;mem[3922] <= 30'b000000000000000000110100110000
                ;mem[3923] <= 30'b000000000000000000110101000000
                ;mem[3924] <= 30'b000000000000000000110101010000
                ;mem[3925] <= 30'b000000000000000000110101100000
                ;mem[3926] <= 30'b000000000000000000110101110000
                ;mem[3927] <= 30'b000000000000000000111011000000
                ;mem[3928] <= 30'b000000000000000000111011010000
                ;mem[3929] <= 30'b000000000000000000111011100000
                ;mem[3930] <= 30'b000000000000000000111011110000
                ;mem[3931] <= 30'b000000000000000000111100000000
                ;mem[3932] <= 30'b000000000000000000111100010000
                ;mem[3933] <= 30'b000000000000000000111100100000
                ;mem[3934] <= 30'b000000000000000000111100110000
                ;mem[3935] <= 30'b000000001000000000000000100000
                ;mem[3936] <= 30'b000000001000000000000000110000
                ;mem[3937] <= 30'b000000001000000000000001000000
                ;mem[3938] <= 30'b000000001000000000000001010000
                ;mem[3939] <= 30'b000000001000000000000001100000
                ;mem[3940] <= 30'b000000001000000000000001110000
                ;mem[3941] <= 30'b000000001000000000000010000000
                ;mem[3942] <= 30'b000000001000000000000010010000
                ;mem[3943] <= 30'b000000001000000000000010100000
                ;mem[3944] <= 30'b000000001000000000000111100000
                ;mem[3945] <= 30'b000000001000000000000111110000
                ;mem[3946] <= 30'b000000001000000000001000000000
                ;mem[3947] <= 30'b000000001000000000001000010000
                ;mem[3948] <= 30'b000000001000000000001000100000
                ;mem[3949] <= 30'b000000001000000000001000110000
                ;mem[3950] <= 30'b000000001000000000001001000000
                ;mem[3951] <= 30'b000000001000000000001001010000
                ;mem[3952] <= 30'b000000001000000000001001100000
                ;mem[3953] <= 30'b000000001000000000001001110000
                ;mem[3954] <= 30'b000000001000000000001111000000
                ;mem[3955] <= 30'b000000001000000000001111010000
                ;mem[3956] <= 30'b000000001000000000001111100000
                ;mem[3957] <= 30'b000000001000000000001111110000
                ;mem[3958] <= 30'b000000001000000000010000000000
                ;mem[3959] <= 30'b000000001000000000010000010000
                ;mem[3960] <= 30'b000000001000000000010000100000
                ;mem[3961] <= 30'b000000001000000000010000110000
                ;mem[3962] <= 30'b000000001000000000010101110000
                ;mem[3963] <= 30'b000000001000000000010110000000
                ;mem[3964] <= 30'b000000001000000000010110010000
                ;mem[3965] <= 30'b000000001000000000010111000000
                ;mem[3966] <= 30'b000000001000000000010111010000
                ;mem[3967] <= 30'b000000001000000000010111100000
                ;mem[3968] <= 30'b000000001000000000010111110000
                ;mem[3969] <= 30'b000000001000000000011000000000
                ;mem[3970] <= 30'b000000001000000000011100100000
                ;mem[3971] <= 30'b000000001000000000011100110000
                ;mem[3972] <= 30'b000000001000000000011101000000
                ;mem[3973] <= 30'b000000001000000000011110010000
                ;mem[3974] <= 30'b000000001000000000011110100000
                ;mem[3975] <= 30'b000000001000000000011110110000
                ;mem[3976] <= 30'b000000001000000000011111000000
                ;mem[3977] <= 30'b000000001000000000100011100000
                ;mem[3978] <= 30'b000000001000000000100011110000
                ;mem[3979] <= 30'b000000001000000000100101100000
                ;mem[3980] <= 30'b000000001000000000100101110000
                ;mem[3981] <= 30'b000000001000000000100110000000
                ;mem[3982] <= 30'b000000001000000000101010100000
                ;mem[3983] <= 30'b000000001000000000101010110000
                ;mem[3984] <= 30'b000000001000000000101100100000
                ;mem[3985] <= 30'b000000001000000000101100110000
                ;mem[3986] <= 30'b000000001000000000101101000000
                ;mem[3987] <= 30'b000000001000000000101101010000
                ;mem[3988] <= 30'b000000001000000000110001010000
                ;mem[3989] <= 30'b000000001000000000110001100000
                ;mem[3990] <= 30'b000000001000000000110011110000
                ;mem[3991] <= 30'b000000001000000000110100000000
                ;mem[3992] <= 30'b000000001000000000110100010000
                ;mem[3993] <= 30'b000000001000000000111000000000
                ;mem[3994] <= 30'b000000001000000000111000010000
                ;mem[3995] <= 30'b000000001000000000111000100000
                ;mem[3996] <= 30'b000000001000000000111010110000
                ;mem[3997] <= 30'b000000001000000000111011000000
                ;mem[3998] <= 30'b000000001000000000111011010000
                ;mem[3999] <= 30'b000000001000000000111111000000
                ;mem[4000] <= 30'b000000001000000000111111010000
                ;mem[4001] <= 30'b000000010000000000000000100000
                ;mem[4002] <= 30'b000000010000000000000000110000
                ;mem[4003] <= 30'b000000010000000000000001000000
                ;mem[4004] <= 30'b000000010000000000000001010000
                ;mem[4005] <= 30'b000000010000000000000101010000
                ;mem[4006] <= 30'b000000010000000000000101100000
                ;mem[4007] <= 30'b000000010000000000000111110000
                ;mem[4008] <= 30'b000000010000000000001000000000
                ;mem[4009] <= 30'b000000010000000000001000010000
                ;mem[4010] <= 30'b000000010000000000001100000000
                ;mem[4011] <= 30'b000000010000000000001100010000
                ;mem[4012] <= 30'b000000010000000000001100100000
                ;mem[4013] <= 30'b000000010000000000001110110000
                ;mem[4014] <= 30'b000000010000000000001111000000
                ;mem[4015] <= 30'b000000010000000000001111010000
                ;mem[4016] <= 30'b000000010000000000010011000000
                ;mem[4017] <= 30'b000000010000000000010011010000
                ;mem[4018] <= 30'b000000010000000000010101110000
                ;mem[4019] <= 30'b000000010000000000010110000000
                ;mem[4020] <= 30'b000000010000000000010110010000
                ;mem[4021] <= 30'b000000010000000000011010000000
                ;mem[4022] <= 30'b000000010000000000011010010000
                ;mem[4023] <= 30'b000000010000000000011100110000
                ;mem[4024] <= 30'b000000010000000000011101000000
                ;mem[4025] <= 30'b000000010000000000011101010000
                ;mem[4026] <= 30'b000000010000000000100001000000
                ;mem[4027] <= 30'b000000010000000000100001010000
                ;mem[4028] <= 30'b000000010000000000100011110000
                ;mem[4029] <= 30'b000000010000000000100100000000
                ;mem[4030] <= 30'b000000010000000000101000000000
                ;mem[4031] <= 30'b000000010000000000101000010000
                ;mem[4032] <= 30'b000000010000000000101000100000
                ;mem[4033] <= 30'b000000010000000000101010110000
                ;mem[4034] <= 30'b000000010000000000101011000000
                ;mem[4035] <= 30'b000000010000000000101111000000
                ;mem[4036] <= 30'b000000010000000000101111010000
                ;mem[4037] <= 30'b000000010000000000101111100000
                ;mem[4038] <= 30'b000000010000000000110001100000
                ;mem[4039] <= 30'b000000010000000000110001110000
                ;mem[4040] <= 30'b000000010000000000110010000000
                ;mem[4041] <= 30'b000000010000000000110110000000
                ;mem[4042] <= 30'b000000010000000000110110010000
                ;mem[4043] <= 30'b000000010000000000110110100000
                ;mem[4044] <= 30'b000000010000000000110110110000
                ;mem[4045] <= 30'b000000010000000000111000010000
                ;mem[4046] <= 30'b000000010000000000111000100000
                ;mem[4047] <= 30'b000000010000000000111000110000
                ;mem[4048] <= 30'b000000010000000000111101000000
                ;mem[4049] <= 30'b000000010000000000111101010000
                ;mem[4050] <= 30'b000000010000000000111101100000
                ;mem[4051] <= 30'b000000010000000000111101110000
                ;mem[4052] <= 30'b000000010000000000111110000000
                ;mem[4053] <= 30'b000000010000000000111110010000
                ;mem[4054] <= 30'b000000010000000000111110100000
                ;mem[4055] <= 30'b000000010000000000111110110000
                ;mem[4056] <= 30'b000000010000000000111111000000
                ;mem[4057] <= 30'b000000010000000000111111010000
                ;mem[4058] <= 30'b000000010000000000111111100000
                ;mem[4059] <= 30'b000000000000000001000011000000
                ;mem[4060] <= 30'b000000000000000001000011010000
                ;mem[4061] <= 30'b000000000000000001000011100000
                ;mem[4062] <= 30'b000000000000000001000101100000
                ;mem[4063] <= 30'b000000000000000001000101110000
                ;mem[4064] <= 30'b000000000000000001000110000000
                ;mem[4065] <= 30'b000000000000000001001010000000
                ;mem[4066] <= 30'b000000000000000001001010010000
                ;mem[4067] <= 30'b000000000000000001001010100000
                ;mem[4068] <= 30'b000000000000000001001010110000
                ;mem[4069] <= 30'b000000000000000001001100010000
                ;mem[4070] <= 30'b000000000000000001001100100000
                ;mem[4071] <= 30'b000000000000000001001100110000
                ;mem[4072] <= 30'b000000000000000001010001000000
                ;mem[4073] <= 30'b000000000000000001010001010000
                ;mem[4074] <= 30'b000000000000000001010001100000
                ;mem[4075] <= 30'b000000000000000001010001110000
                ;mem[4076] <= 30'b000000000000000001010010000000
                ;mem[4077] <= 30'b000000000000000001010010010000
                ;mem[4078] <= 30'b000000000000000001010010100000
                ;mem[4079] <= 30'b000000000000000001010010110000
                ;mem[4080] <= 30'b000000000000000001010011000000
                ;mem[4081] <= 30'b000000000000000001010011010000
                ;mem[4082] <= 30'b000000000000000001010011100000
                ;mem[4083] <= 30'b000000000000000001011000010000
                ;mem[4084] <= 30'b000000000000000001011000100000
                ;mem[4085] <= 30'b000000000000000001011000110000
                ;mem[4086] <= 30'b000000000000000001011001000000
                ;mem[4087] <= 30'b000000000000000001011001010000
                ;mem[4088] <= 30'b000000000000000001011001100000
                ;mem[4089] <= 30'b000000000000000001011001110000
                ;mem[4090] <= 30'b000000000000000001011010000000
                ;mem[4091] <= 30'b000000000000000001011010010000
                ;mem[4092] <= 30'b000000000000000001011111100000
                ;mem[4093] <= 30'b000000000000000001011111110000
                ;mem[4094] <= 30'b000000000000000001100000000000
                ;mem[4095] <= 30'b000000000000000001100000010000
                ;mem[4096] <= 30'b000000000000000001100000100000
                ;mem[4097] <= 30'b000000000000000001100000110000
                ;mem[4098] <= 30'b000000000000000001100001000000
                ;mem[4099] <= 30'b000000000000000001100111000000
                ;mem[4100] <= 30'b000000000000000001100111010000
                ;mem[4101] <= 30'b000000000000000000011110110000
                ;mem[4102] <= 30'b000000000000000000011111000000
                ;mem[4103] <= 30'b000000000000000000100101110000
                ;mem[4104] <= 30'b000000000000000000100110000000
                ;mem[4105] <= 30'b000000000000000000101100110000
                ;mem[4106] <= 30'b000000000000000000101101000000
                ;mem[4107] <= 30'b000000000000000000101101010000
                ;mem[4108] <= 30'b000000000000000000110100000000
                ;mem[4109] <= 30'b000000000000000000110100010000
                ;mem[4110] <= 30'b000000000000000000111011010000
                ;mem[4111] <= 30'b000000000000000000111011100000
                ;mem[4112] <= 30'b000000001000000000000000110000
                ;mem[4113] <= 30'b000000001000000000000001000000
                ;mem[4114] <= 30'b000000001000000000000001010000
                ;mem[4115] <= 30'b000000001000000000001000000000
                ;mem[4116] <= 30'b000000001000000000001000010000
                ;mem[4117] <= 30'b000000001000000000001111010000
                ;mem[4118] <= 30'b000000001000000000001111100000
                ;mem[4119] <= 30'b000000001000000000010110010000
                ;mem[4120] <= 30'b000000001000000000010110100000
                ;mem[4121] <= 30'b000000001000000000011101000000
                ;mem[4122] <= 30'b000000001000000000011101010000
                ;mem[4123] <= 30'b000000001000000000011101100000
                ;mem[4124] <= 30'b000000001000000000100100010000
                ;mem[4125] <= 30'b000000001000000000100100100000
                ;mem[4126] <= 30'b000000001000000000101011000000
                ;mem[4127] <= 30'b000000001000000000101011010000
                ;mem[4128] <= 30'b000000001000000000101011100000
                ;mem[4129] <= 30'b000000001000000000110010000000
                ;mem[4130] <= 30'b000000001000000000110010010000
                ;mem[4131] <= 30'b000000001000000000110010100000
                ;mem[4132] <= 30'b000000001000000000111001010000
                ;mem[4133] <= 30'b000000001000000000111001100000
                ;mem[4134] <= 30'b000000001000000000111001110000
                ;mem[4135] <= 30'b000000010000000000000110000000
                ;mem[4136] <= 30'b000000010000000000000110010000
                ;mem[4137] <= 30'b000000010000000000000110100000
                ;mem[4138] <= 30'b000000010000000000001101010000
                ;mem[4139] <= 30'b000000010000000000001101100000
                ;mem[4140] <= 30'b000000010000000000001101110000
                ;mem[4141] <= 30'b000000010000000000010100100000
                ;mem[4142] <= 30'b000000010000000000010100110000
                ;mem[4143] <= 30'b000000010000000000011011100000
                ;mem[4144] <= 30'b000000010000000000011011110000
                ;mem[4145] <= 30'b000000010000000000100010100000
                ;mem[4146] <= 30'b000000010000000000100010110000
                ;mem[4147] <= 30'b000000010000000000101001100000
                ;mem[4148] <= 30'b000000010000000000101001110000
                ;mem[4149] <= 30'b000000010000000000110000010000
                ;mem[4150] <= 30'b000000010000000000110000100000
                ;mem[4151] <= 30'b000000010000000000110000110000
                ;mem[4152] <= 30'b000000010000000000110111010000
                ;mem[4153] <= 30'b000000010000000000110111100000
                ;mem[4154] <= 30'b000000010000000000110111110000
                ;mem[4155] <= 30'b000000010000000000111110100000
                ;mem[4156] <= 30'b000000010000000000111110110000
                ;mem[4157] <= 30'b000000000000000001000100010000
                ;mem[4158] <= 30'b000000000000000001000100100000
                ;mem[4159] <= 30'b000000000000000001000100110000
                ;mem[4160] <= 30'b000000000000000001001011010000
                ;mem[4161] <= 30'b000000000000000001001011100000
                ;mem[4162] <= 30'b000000000000000001001011110000
                ;mem[4163] <= 30'b000000000000000001010010100000
                ;mem[4164] <= 30'b000000000000000001010010110000
                ;mem[4165] <= 30'b000000000000000001011001100000
                ;mem[4166] <= 30'b000000000000000001011001110000
                ;mem[4167] <= 30'b000000000000000001100000100000
                ;mem[4168] <= 30'b000000000000000001100000110000
                ;mem[4169] <= 30'b000000000000000000101100010000
                ;mem[4170] <= 30'b000000000000000000101100100000
                ;mem[4171] <= 30'b000000000000000000101100110000
                ;mem[4172] <= 30'b000000000000000000101101000000
                ;mem[4173] <= 30'b000000000000000000101101010000
                ;mem[4174] <= 30'b000000000000000000101101100000
                ;mem[4175] <= 30'b000000000000000000101101110000
                ;mem[4176] <= 30'b000000000000000000110010110000
                ;mem[4177] <= 30'b000000000000000000110011000000
                ;mem[4178] <= 30'b000000000000000000110011010000
                ;mem[4179] <= 30'b000000000000000000110011100000
                ;mem[4180] <= 30'b000000000000000000110011110000
                ;mem[4181] <= 30'b000000000000000000110100000000
                ;mem[4182] <= 30'b000000000000000000110100010000
                ;mem[4183] <= 30'b000000000000000000110100100000
                ;mem[4184] <= 30'b000000000000000000110100110000
                ;mem[4185] <= 30'b000000000000000000110101000000
                ;mem[4186] <= 30'b000000000000000000111001110000
                ;mem[4187] <= 30'b000000000000000000111010000000
                ;mem[4188] <= 30'b000000000000000000111010010000
                ;mem[4189] <= 30'b000000000000000000111010100000
                ;mem[4190] <= 30'b000000000000000000111011000000
                ;mem[4191] <= 30'b000000000000000000111011010000
                ;mem[4192] <= 30'b000000000000000000111011100000
                ;mem[4193] <= 30'b000000000000000000111011110000
                ;mem[4194] <= 30'b000000000000000000111100000000
                ;mem[4195] <= 30'b000000000000000000111100010000
                ;mem[4196] <= 30'b000000001000000000000000010000
                ;mem[4197] <= 30'b000000001000000000000000100000
                ;mem[4198] <= 30'b000000001000000000000000110000
                ;mem[4199] <= 30'b000000001000000000000001000000
                ;mem[4200] <= 30'b000000001000000000000001010000
                ;mem[4201] <= 30'b000000001000000000000001100000
                ;mem[4202] <= 30'b000000001000000000000001110000
                ;mem[4203] <= 30'b000000001000000000000110110000
                ;mem[4204] <= 30'b000000001000000000000111000000
                ;mem[4205] <= 30'b000000001000000000000111010000
                ;mem[4206] <= 30'b000000001000000000000111100000
                ;mem[4207] <= 30'b000000001000000000000111110000
                ;mem[4208] <= 30'b000000001000000000001000000000
                ;mem[4209] <= 30'b000000001000000000001000010000
                ;mem[4210] <= 30'b000000001000000000001000100000
                ;mem[4211] <= 30'b000000001000000000001000110000
                ;mem[4212] <= 30'b000000001000000000001001000000
                ;mem[4213] <= 30'b000000001000000000001101110000
                ;mem[4214] <= 30'b000000001000000000001110000000
                ;mem[4215] <= 30'b000000001000000000001110010000
                ;mem[4216] <= 30'b000000001000000000001110100000
                ;mem[4217] <= 30'b000000001000000000001111000000
                ;mem[4218] <= 30'b000000001000000000001111010000
                ;mem[4219] <= 30'b000000001000000000001111100000
                ;mem[4220] <= 30'b000000001000000000001111110000
                ;mem[4221] <= 30'b000000001000000000010000000000
                ;mem[4222] <= 30'b000000001000000000010000010000
                ;mem[4223] <= 30'b000000001000000000010101000000
                ;mem[4224] <= 30'b000000001000000000010110100000
                ;mem[4225] <= 30'b000000001000000000010110110000
                ;mem[4226] <= 30'b000000001000000000010111000000
                ;mem[4227] <= 30'b000000001000000000011101010000
                ;mem[4228] <= 30'b000000001000000000011101100000
                ;mem[4229] <= 30'b000000001000000000011101110000
                ;mem[4230] <= 30'b000000001000000000011110000000
                ;mem[4231] <= 30'b000000001000000000100100000000
                ;mem[4232] <= 30'b000000001000000000100100010000
                ;mem[4233] <= 30'b000000001000000000100100100000
                ;mem[4234] <= 30'b000000001000000000100100110000
                ;mem[4235] <= 30'b000000001000000000101010110000
                ;mem[4236] <= 30'b000000001000000000101011000000
                ;mem[4237] <= 30'b000000001000000000101011010000
                ;mem[4238] <= 30'b000000001000000000101011100000
                ;mem[4239] <= 30'b000000001000000000101011110000
                ;mem[4240] <= 30'b000000001000000000110001110000
                ;mem[4241] <= 30'b000000001000000000110010000000
                ;mem[4242] <= 30'b000000001000000000110010010000
                ;mem[4243] <= 30'b000000001000000000110010100000
                ;mem[4244] <= 30'b000000001000000000110010110000
                ;mem[4245] <= 30'b000000001000000000110011000000
                ;mem[4246] <= 30'b000000001000000000111001010000
                ;mem[4247] <= 30'b000000001000000000111001100000
                ;mem[4248] <= 30'b000000001000000000111001110000
                ;mem[4249] <= 30'b000000001000000000111010000000
                ;mem[4250] <= 30'b000000001000000000111010010000
                ;mem[4251] <= 30'b000000001000000000111010100000
                ;mem[4252] <= 30'b000000010000000000000101110000
                ;mem[4253] <= 30'b000000010000000000000110000000
                ;mem[4254] <= 30'b000000010000000000000110010000
                ;mem[4255] <= 30'b000000010000000000000110100000
                ;mem[4256] <= 30'b000000010000000000000110110000
                ;mem[4257] <= 30'b000000010000000000000111000000
                ;mem[4258] <= 30'b000000010000000000001101010000
                ;mem[4259] <= 30'b000000010000000000001101100000
                ;mem[4260] <= 30'b000000010000000000001101110000
                ;mem[4261] <= 30'b000000010000000000001110000000
                ;mem[4262] <= 30'b000000010000000000001110010000
                ;mem[4263] <= 30'b000000010000000000001110100000
                ;mem[4264] <= 30'b000000010000000000010100110000
                ;mem[4265] <= 30'b000000010000000000010101000000
                ;mem[4266] <= 30'b000000010000000000010101010000
                ;mem[4267] <= 30'b000000010000000000010101100000
                ;mem[4268] <= 30'b000000010000000000010101110000
                ;mem[4269] <= 30'b000000010000000000011100010000
                ;mem[4270] <= 30'b000000010000000000011100100000
                ;mem[4271] <= 30'b000000010000000000011100110000
                ;mem[4272] <= 30'b000000010000000000100011010000
                ;mem[4273] <= 30'b000000010000000000100011100000
                ;mem[4274] <= 30'b000000010000000000100011110000
                ;mem[4275] <= 30'b000000010000000000101010000000
                ;mem[4276] <= 30'b000000010000000000101010010000
                ;mem[4277] <= 30'b000000010000000000101010100000
                ;mem[4278] <= 30'b000000010000000000110000110000
                ;mem[4279] <= 30'b000000010000000000110001000000
                ;mem[4280] <= 30'b000000010000000000110001010000
                ;mem[4281] <= 30'b000000010000000000110001100000
                ;mem[4282] <= 30'b000000010000000000110111100000
                ;mem[4283] <= 30'b000000010000000000110111110000
                ;mem[4284] <= 30'b000000010000000000111000000000
                ;mem[4285] <= 30'b000000010000000000111000010000
                ;mem[4286] <= 30'b000000010000000000111110000000
                ;mem[4287] <= 30'b000000010000000000111110010000
                ;mem[4288] <= 30'b000000010000000000111110100000
                ;mem[4289] <= 30'b000000010000000000111110110000
                ;mem[4290] <= 30'b000000010000000000111111000000
                ;mem[4291] <= 30'b000000000000000001000100110000
                ;mem[4292] <= 30'b000000000000000001000101000000
                ;mem[4293] <= 30'b000000000000000001000101010000
                ;mem[4294] <= 30'b000000000000000001000101100000
                ;mem[4295] <= 30'b000000000000000001001011100000
                ;mem[4296] <= 30'b000000000000000001001011110000
                ;mem[4297] <= 30'b000000000000000001001100000000
                ;mem[4298] <= 30'b000000000000000001001100010000
                ;mem[4299] <= 30'b000000000000000001010010000000
                ;mem[4300] <= 30'b000000000000000001010010010000
                ;mem[4301] <= 30'b000000000000000001010010100000
                ;mem[4302] <= 30'b000000000000000001010010110000
                ;mem[4303] <= 30'b000000000000000001010011000000
                ;mem[4304] <= 30'b000000000000000001011000010000
                ;mem[4305] <= 30'b000000000000000001011000100000
                ;mem[4306] <= 30'b000000000000000001011000110000
                ;mem[4307] <= 30'b000000000000000001011001000000
                ;mem[4308] <= 30'b000000000000000001011001010000
                ;mem[4309] <= 30'b000000000000000001011001100000
                ;mem[4310] <= 30'b000000000000000001011111000000
                ;mem[4311] <= 30'b000000000000000001011111010000
                ;mem[4312] <= 30'b000000000000000001011111100000
                ;mem[4313] <= 30'b000000000000000001011111110000
                ;mem[4314] <= 30'b000000000000000001100000000000
                ;mem[4315] <= 30'b000000000000000001100000010000
                ;mem[4316] <= 30'b000000000000000001100110000000
                ;mem[4317] <= 30'b000000000000000001100110010000
                ;mem[4318] <= 30'b000000000000000001100110100000
                ;mem[4319] <= 30'b000000000000000001100110110000
                ;mem[4320] <= 30'b000000000000000001101101010000
                ;mem[4321] <= 30'b000000000000000000100110000000
                ;mem[4322] <= 30'b000000000000000000100110010000
                ;mem[4323] <= 30'b000000000000000000101101000000
                ;mem[4324] <= 30'b000000000000000000101101010000
                ;mem[4325] <= 30'b000000000000000000101101100000
                ;mem[4326] <= 30'b000000000000000000110100010000
                ;mem[4327] <= 30'b000000000000000000110100100000
                ;mem[4328] <= 30'b000000000000000000111011010000
                ;mem[4329] <= 30'b000000000000000000111011100000
                ;mem[4330] <= 30'b000000001000000000000001000000
                ;mem[4331] <= 30'b000000001000000000000001010000
                ;mem[4332] <= 30'b000000001000000000000001100000
                ;mem[4333] <= 30'b000000001000000000001000010000
                ;mem[4334] <= 30'b000000001000000000001000100000
                ;mem[4335] <= 30'b000000001000000000001111010000
                ;mem[4336] <= 30'b000000001000000000001111100000
                ;mem[4337] <= 30'b000000001000000000010110010000
                ;mem[4338] <= 30'b000000001000000000010110100000
                ;mem[4339] <= 30'b000000001000000000011101010000
                ;mem[4340] <= 30'b000000001000000000011101100000
                ;mem[4341] <= 30'b000000001000000000100100010000
                ;mem[4342] <= 30'b000000001000000000100100100000
                ;mem[4343] <= 30'b000000001000000000100100110000
                ;mem[4344] <= 30'b000000001000000000101011010000
                ;mem[4345] <= 30'b000000001000000000101011100000
                ;mem[4346] <= 30'b000000001000000000101011110000
                ;mem[4347] <= 30'b000000001000000000110010100000
                ;mem[4348] <= 30'b000000001000000000110010110000
                ;mem[4349] <= 30'b000000001000000000111001100000
                ;mem[4350] <= 30'b000000001000000000111001110000
                ;mem[4351] <= 30'b000000010000000000000110100000
                ;mem[4352] <= 30'b000000010000000000000110110000
                ;mem[4353] <= 30'b000000010000000000001101100000
                ;mem[4354] <= 30'b000000010000000000001101110000
                ;mem[4355] <= 30'b000000010000000000010100100000
                ;mem[4356] <= 30'b000000010000000000010100110000
                ;mem[4357] <= 30'b000000010000000000011011100000
                ;mem[4358] <= 30'b000000010000000000011011110000
                ;mem[4359] <= 30'b000000010000000000011100000000
                ;mem[4360] <= 30'b000000010000000000100010110000
                ;mem[4361] <= 30'b000000010000000000100011000000
                ;mem[4362] <= 30'b000000010000000000101001110000
                ;mem[4363] <= 30'b000000010000000000101010000000
                ;mem[4364] <= 30'b000000010000000000110000110000
                ;mem[4365] <= 30'b000000010000000000110001000000
                ;mem[4366] <= 30'b000000010000000000110111110000
                ;mem[4367] <= 30'b000000010000000000111000000000
                ;mem[4368] <= 30'b000000010000000000111110110000
                ;mem[4369] <= 30'b000000010000000000111111000000
                ;mem[4370] <= 30'b000000000000000001000100110000
                ;mem[4371] <= 30'b000000000000000001000101000000
                ;mem[4372] <= 30'b000000000000000001001011110000
                ;mem[4373] <= 30'b000000000000000001001100000000
                ;mem[4374] <= 30'b000000000000000001010010110000
                ;mem[4375] <= 30'b000000000000000001010011000000
                ;mem[4376] <= 30'b000000000000000001011001110000
                ;mem[4377] <= 30'b000000000000000001011010000000
                ;mem[4378] <= 30'b000000000000000001100000110000
                ;mem[4379] <= 30'b000000000000000001100001000000
                ;mem[4380] <= 30'b000000000000000001101000000000
                ;mem[4381] <= 30'b000000000000000000100101010000
                ;mem[4382] <= 30'b000000000000000000100101100000
                ;mem[4383] <= 30'b000000000000000000100101110000
                ;mem[4384] <= 30'b000000000000000000100110000000
                ;mem[4385] <= 30'b000000000000000000100110010000
                ;mem[4386] <= 30'b000000000000000000101011110000
                ;mem[4387] <= 30'b000000000000000000101100000000
                ;mem[4388] <= 30'b000000000000000000101100010000
                ;mem[4389] <= 30'b000000000000000000101100100000
                ;mem[4390] <= 30'b000000000000000000101100110000
                ;mem[4391] <= 30'b000000000000000000101101000000
                ;mem[4392] <= 30'b000000000000000000101101010000
                ;mem[4393] <= 30'b000000000000000000101101100000
                ;mem[4394] <= 30'b000000000000000000101101110000
                ;mem[4395] <= 30'b000000000000000000110010110000
                ;mem[4396] <= 30'b000000000000000000110011000000
                ;mem[4397] <= 30'b000000000000000000110011010000
                ;mem[4398] <= 30'b000000000000000000110011100000
                ;mem[4399] <= 30'b000000000000000000110011110000
                ;mem[4400] <= 30'b000000000000000000110100100000
                ;mem[4401] <= 30'b000000000000000000110100110000
                ;mem[4402] <= 30'b000000000000000000111001110000
                ;mem[4403] <= 30'b000000000000000000111010000000
                ;mem[4404] <= 30'b000000000000000000111011100000
                ;mem[4405] <= 30'b000000000000000000111011110000
                ;mem[4406] <= 30'b000000001000000000000000000000
                ;mem[4407] <= 30'b000000001000000000000000010000
                ;mem[4408] <= 30'b000000001000000000000000100000
                ;mem[4409] <= 30'b000000001000000000000000110000
                ;mem[4410] <= 30'b000000001000000000000001000000
                ;mem[4411] <= 30'b000000001000000000000001010000
                ;mem[4412] <= 30'b000000001000000000000001100000
                ;mem[4413] <= 30'b000000001000000000000001110000
                ;mem[4414] <= 30'b000000001000000000000110110000
                ;mem[4415] <= 30'b000000001000000000000111000000
                ;mem[4416] <= 30'b000000001000000000000111010000
                ;mem[4417] <= 30'b000000001000000000000111100000
                ;mem[4418] <= 30'b000000001000000000000111110000
                ;mem[4419] <= 30'b000000001000000000001000100000
                ;mem[4420] <= 30'b000000001000000000001000110000
                ;mem[4421] <= 30'b000000001000000000001101110000
                ;mem[4422] <= 30'b000000001000000000001110000000
                ;mem[4423] <= 30'b000000001000000000001111100000
                ;mem[4424] <= 30'b000000001000000000001111110000
                ;mem[4425] <= 30'b000000001000000000010110100000
                ;mem[4426] <= 30'b000000001000000000010110110000
                ;mem[4427] <= 30'b000000001000000000011101010000
                ;mem[4428] <= 30'b000000001000000000011101100000
                ;mem[4429] <= 30'b000000001000000000011101110000
                ;mem[4430] <= 30'b000000001000000000100100000000
                ;mem[4431] <= 30'b000000001000000000100100010000
                ;mem[4432] <= 30'b000000001000000000100100100000
                ;mem[4433] <= 30'b000000001000000000101010110000
                ;mem[4434] <= 30'b000000001000000000101011000000
                ;mem[4435] <= 30'b000000001000000000101011010000
                ;mem[4436] <= 30'b000000001000000000101011100000
                ;mem[4437] <= 30'b000000001000000000110001010000
                ;mem[4438] <= 30'b000000001000000000110001100000
                ;mem[4439] <= 30'b000000001000000000110001110000
                ;mem[4440] <= 30'b000000001000000000110010000000
                ;mem[4441] <= 30'b000000001000000000110010010000
                ;mem[4442] <= 30'b000000001000000000110010100000
                ;mem[4443] <= 30'b000000001000000000110010110000
                ;mem[4444] <= 30'b000000001000000000111000010000
                ;mem[4445] <= 30'b000000001000000000111000100000
                ;mem[4446] <= 30'b000000001000000000111000110000
                ;mem[4447] <= 30'b000000001000000000111001000000
                ;mem[4448] <= 30'b000000001000000000111001010000
                ;mem[4449] <= 30'b000000001000000000111001100000
                ;mem[4450] <= 30'b000000001000000000111001110000
                ;mem[4451] <= 30'b000000001000000000111010000000
                ;mem[4452] <= 30'b000000001000000000111010010000
                ;mem[4453] <= 30'b000000001000000000111111010000
                ;mem[4454] <= 30'b000000001000000000111111100000
                ;mem[4455] <= 30'b000000001000000000111111110000
                ;mem[4456] <= 30'b000000010000000000000101010000
                ;mem[4457] <= 30'b000000010000000000000101100000
                ;mem[4458] <= 30'b000000010000000000000101110000
                ;mem[4459] <= 30'b000000010000000000000110000000
                ;mem[4460] <= 30'b000000010000000000000110010000
                ;mem[4461] <= 30'b000000010000000000000110100000
                ;mem[4462] <= 30'b000000010000000000000110110000
                ;mem[4463] <= 30'b000000010000000000001100010000
                ;mem[4464] <= 30'b000000010000000000001100100000
                ;mem[4465] <= 30'b000000010000000000001100110000
                ;mem[4466] <= 30'b000000010000000000001101000000
                ;mem[4467] <= 30'b000000010000000000001101010000
                ;mem[4468] <= 30'b000000010000000000001101100000
                ;mem[4469] <= 30'b000000010000000000001101110000
                ;mem[4470] <= 30'b000000010000000000001110000000
                ;mem[4471] <= 30'b000000010000000000001110010000
                ;mem[4472] <= 30'b000000010000000000010011010000
                ;mem[4473] <= 30'b000000010000000000010011100000
                ;mem[4474] <= 30'b000000010000000000010011110000
                ;mem[4475] <= 30'b000000010000000000010100110000
                ;mem[4476] <= 30'b000000010000000000010101000000
                ;mem[4477] <= 30'b000000010000000000010101010000
                ;mem[4478] <= 30'b000000010000000000010101100000
                ;mem[4479] <= 30'b000000010000000000011100000000
                ;mem[4480] <= 30'b000000010000000000011100010000
                ;mem[4481] <= 30'b000000010000000000011100100000
                ;mem[4482] <= 30'b000000010000000000011100110000
                ;mem[4483] <= 30'b000000010000000000100011010000
                ;mem[4484] <= 30'b000000010000000000100011100000
                ;mem[4485] <= 30'b000000010000000000100011110000
                ;mem[4486] <= 30'b000000010000000000101010100000
                ;mem[4487] <= 30'b000000010000000000101010110000
                ;mem[4488] <= 30'b000000010000000000101011000000
                ;mem[4489] <= 30'b000000010000000000110001110000
                ;mem[4490] <= 30'b000000010000000000110010000000
                ;mem[4491] <= 30'b000000010000000000111000100000
                ;mem[4492] <= 30'b000000010000000000111000110000
                ;mem[4493] <= 30'b000000010000000000111001000000
                ;mem[4494] <= 30'b000000010000000000111111000000
                ;mem[4495] <= 30'b000000010000000000111111010000
                ;mem[4496] <= 30'b000000010000000000111111100000
                ;mem[4497] <= 30'b000000010000000000111111110000
                ;mem[4498] <= 30'b000000000000000001000101110000
                ;mem[4499] <= 30'b000000000000000001000110000000
                ;mem[4500] <= 30'b000000000000000001001100100000
                ;mem[4501] <= 30'b000000000000000001001100110000
                ;mem[4502] <= 30'b000000000000000001001101000000
                ;mem[4503] <= 30'b000000000000000001010011000000
                ;mem[4504] <= 30'b000000000000000001010011010000
                ;mem[4505] <= 30'b000000000000000001010011100000
                ;mem[4506] <= 30'b000000000000000001010011110000
                ;mem[4507] <= 30'b000000000000000001010100000000
                ;mem[4508] <= 30'b000000000000000001011001010000
                ;mem[4509] <= 30'b000000000000000001011001100000
                ;mem[4510] <= 30'b000000000000000001011001110000
                ;mem[4511] <= 30'b000000000000000001011010000000
                ;mem[4512] <= 30'b000000000000000001011010010000
                ;mem[4513] <= 30'b000000000000000001011010100000
                ;mem[4514] <= 30'b000000000000000001011010110000
                ;mem[4515] <= 30'b000000000000000001011111100000
                ;mem[4516] <= 30'b000000000000000001011111110000
                ;mem[4517] <= 30'b000000000000000001100000000000
                ;mem[4518] <= 30'b000000000000000001100000010000
                ;mem[4519] <= 30'b000000000000000001100000100000
                ;mem[4520] <= 30'b000000000000000001100000110000
                ;mem[4521] <= 30'b000000000000000001100001000000
                ;mem[4522] <= 30'b000000000000000001100001010000
                ;mem[4523] <= 30'b000000000000000001100110100000
                ;mem[4524] <= 30'b000000000000000001100110110000
                ;mem[4525] <= 30'b000000000000000001100111000000
                ;mem[4526] <= 30'b000000000000000001100111010000
                ;mem[4527] <= 30'b000000000000000001100111100000
                ;mem[4528] <= 30'b000000000000000000100101100000
                ;mem[4529] <= 30'b000000000000000000100101110000
                ;mem[4530] <= 30'b000000000000000000101100100000
                ;mem[4531] <= 30'b000000000000000000101100110000
                ;mem[4532] <= 30'b000000000000000000101111110000
                ;mem[4533] <= 30'b000000000000000000110000000000
                ;mem[4534] <= 30'b000000000000000000110011110000
                ;mem[4535] <= 30'b000000000000000000110110110000
                ;mem[4536] <= 30'b000000000000000000110111000000
                ;mem[4537] <= 30'b000000000000000000111010100000
                ;mem[4538] <= 30'b000000000000000000111010110000
                ;mem[4539] <= 30'b000000000000000000111101100000
                ;mem[4540] <= 30'b000000000000000000111101110000
                ;mem[4541] <= 30'b000000000000000000111110000000
                ;mem[4542] <= 30'b000000001000000000000000100000
                ;mem[4543] <= 30'b000000001000000000000000110000
                ;mem[4544] <= 30'b000000001000000000000011110000
                ;mem[4545] <= 30'b000000001000000000000100000000
                ;mem[4546] <= 30'b000000001000000000000111110000
                ;mem[4547] <= 30'b000000001000000000001010110000
                ;mem[4548] <= 30'b000000001000000000001011000000
                ;mem[4549] <= 30'b000000001000000000001110100000
                ;mem[4550] <= 30'b000000001000000000001110110000
                ;mem[4551] <= 30'b000000001000000000010001100000
                ;mem[4552] <= 30'b000000001000000000010001110000
                ;mem[4553] <= 30'b000000001000000000010010000000
                ;mem[4554] <= 30'b000000001000000000010101100000
                ;mem[4555] <= 30'b000000001000000000010101110000
                ;mem[4556] <= 30'b000000001000000000011000100000
                ;mem[4557] <= 30'b000000001000000000011000110000
                ;mem[4558] <= 30'b000000001000000000011100100000
                ;mem[4559] <= 30'b000000001000000000011100110000
                ;mem[4560] <= 30'b000000001000000000011111100000
                ;mem[4561] <= 30'b000000001000000000011111110000
                ;mem[4562] <= 30'b000000001000000000100011010000
                ;mem[4563] <= 30'b000000001000000000100011100000
                ;mem[4564] <= 30'b000000001000000000100011110000
                ;mem[4565] <= 30'b000000001000000000100110100000
                ;mem[4566] <= 30'b000000001000000000100110110000
                ;mem[4567] <= 30'b000000001000000000101010000000
                ;mem[4568] <= 30'b000000001000000000101010010000
                ;mem[4569] <= 30'b000000001000000000101010100000
                ;mem[4570] <= 30'b000000001000000000101101010000
                ;mem[4571] <= 30'b000000001000000000101101100000
                ;mem[4572] <= 30'b000000001000000000101101110000
                ;mem[4573] <= 30'b000000001000000000110001000000
                ;mem[4574] <= 30'b000000001000000000110001010000
                ;mem[4575] <= 30'b000000001000000000110001100000
                ;mem[4576] <= 30'b000000001000000000110100010000
                ;mem[4577] <= 30'b000000001000000000110100100000
                ;mem[4578] <= 30'b000000001000000000110100110000
                ;mem[4579] <= 30'b000000001000000000110111110000
                ;mem[4580] <= 30'b000000001000000000111000000000
                ;mem[4581] <= 30'b000000001000000000111000010000
                ;mem[4582] <= 30'b000000001000000000111011010000
                ;mem[4583] <= 30'b000000001000000000111011100000
                ;mem[4584] <= 30'b000000001000000000111110110000
                ;mem[4585] <= 30'b000000001000000000111111000000
                ;mem[4586] <= 30'b000000001000000000111111010000
                ;mem[4587] <= 30'b000000010000000000000001010000
                ;mem[4588] <= 30'b000000010000000000000001100000
                ;mem[4589] <= 30'b000000010000000000000001110000
                ;mem[4590] <= 30'b000000010000000000000101000000
                ;mem[4591] <= 30'b000000010000000000000101010000
                ;mem[4592] <= 30'b000000010000000000000101100000
                ;mem[4593] <= 30'b000000010000000000001000010000
                ;mem[4594] <= 30'b000000010000000000001000100000
                ;mem[4595] <= 30'b000000010000000000001000110000
                ;mem[4596] <= 30'b000000010000000000001011110000
                ;mem[4597] <= 30'b000000010000000000001100000000
                ;mem[4598] <= 30'b000000010000000000001100010000
                ;mem[4599] <= 30'b000000010000000000001111010000
                ;mem[4600] <= 30'b000000010000000000001111100000
                ;mem[4601] <= 30'b000000010000000000010010110000
                ;mem[4602] <= 30'b000000010000000000010011000000
                ;mem[4603] <= 30'b000000010000000000010011010000
                ;mem[4604] <= 30'b000000010000000000010110010000
                ;mem[4605] <= 30'b000000010000000000010110100000
                ;mem[4606] <= 30'b000000010000000000011001100000
                ;mem[4607] <= 30'b000000010000000000011001110000
                ;mem[4608] <= 30'b000000010000000000011010000000
                ;mem[4609] <= 30'b000000010000000000011101010000
                ;mem[4610] <= 30'b000000010000000000011101100000
                ;mem[4611] <= 30'b000000010000000000100000010000
                ;mem[4612] <= 30'b000000010000000000100000100000
                ;mem[4613] <= 30'b000000010000000000100000110000
                ;mem[4614] <= 30'b000000010000000000100001000000
                ;mem[4615] <= 30'b000000010000000000100001010000
                ;mem[4616] <= 30'b000000010000000000100001100000
                ;mem[4617] <= 30'b000000010000000000100001110000
                ;mem[4618] <= 30'b000000010000000000100010000000
                ;mem[4619] <= 30'b000000010000000000100010010000
                ;mem[4620] <= 30'b000000010000000000100010100000
                ;mem[4621] <= 30'b000000010000000000100010110000
                ;mem[4622] <= 30'b000000010000000000100011000000
                ;mem[4623] <= 30'b000000010000000000100011010000
                ;mem[4624] <= 30'b000000010000000000100100010000
                ;mem[4625] <= 30'b000000010000000000100100100000
                ;mem[4626] <= 30'b000000010000000000100111010000
                ;mem[4627] <= 30'b000000010000000000100111100000
                ;mem[4628] <= 30'b000000010000000000100111110000
                ;mem[4629] <= 30'b000000010000000000101000000000
                ;mem[4630] <= 30'b000000010000000000101000010000
                ;mem[4631] <= 30'b000000010000000000101000100000
                ;mem[4632] <= 30'b000000010000000000101000110000
                ;mem[4633] <= 30'b000000010000000000101001000000
                ;mem[4634] <= 30'b000000010000000000101001010000
                ;mem[4635] <= 30'b000000010000000000101001100000
                ;mem[4636] <= 30'b000000010000000000101001110000
                ;mem[4637] <= 30'b000000010000000000101010000000
                ;mem[4638] <= 30'b000000010000000000101010010000
                ;mem[4639] <= 30'b000000010000000000101010100000
                ;mem[4640] <= 30'b000000010000000000101010110000
                ;mem[4641] <= 30'b000000010000000000101011000000
                ;mem[4642] <= 30'b000000010000000000101011010000
                ;mem[4643] <= 30'b000000010000000000101110100000
                ;mem[4644] <= 30'b000000010000000000101110110000
                ;mem[4645] <= 30'b000000010000000000101111000000
                ;mem[4646] <= 30'b000000010000000000101111010000
                ;mem[4647] <= 30'b000000010000000000101111100000
                ;mem[4648] <= 30'b000000010000000000101111110000
                ;mem[4649] <= 30'b000000010000000000110001110000
                ;mem[4650] <= 30'b000000010000000000110010000000
                ;mem[4651] <= 30'b000000010000000000110010010000
                ;mem[4652] <= 30'b000000010000000000111000110000
                ;mem[4653] <= 30'b000000010000000000111001000000
                ;mem[4654] <= 30'b000000010000000000111001010000
                ;mem[4655] <= 30'b000000000000000001000010100000
                ;mem[4656] <= 30'b000000000000000001000010110000
                ;mem[4657] <= 30'b000000000000000001000011000000
                ;mem[4658] <= 30'b000000000000000001000011010000
                ;mem[4659] <= 30'b000000000000000001000011100000
                ;mem[4660] <= 30'b000000000000000001000011110000
                ;mem[4661] <= 30'b000000000000000001000101110000
                ;mem[4662] <= 30'b000000000000000001000110000000
                ;mem[4663] <= 30'b000000000000000001000110010000
                ;mem[4664] <= 30'b000000000000000001001100110000
                ;mem[4665] <= 30'b000000000000000001001101000000
                ;mem[4666] <= 30'b000000000000000001001101010000
                ;mem[4667] <= 30'b000000000000000000101011110000
                ;mem[4668] <= 30'b000000000000000000101100000000
                ;mem[4669] <= 30'b000000000000000000101110110000
                ;mem[4670] <= 30'b000000000000000000101111000000
                ;mem[4671] <= 30'b000000000000000000101111010000
                ;mem[4672] <= 30'b000000000000000000110011000000
                ;mem[4673] <= 30'b000000000000000000110011010000
                ;mem[4674] <= 30'b000000000000000000110011100000
                ;mem[4675] <= 30'b000000000000000000110011110000
                ;mem[4676] <= 30'b000000000000000000110100000000
                ;mem[4677] <= 30'b000000000000000000110100010000
                ;mem[4678] <= 30'b000000000000000000110100100000
                ;mem[4679] <= 30'b000000000000000000110100110000
                ;mem[4680] <= 30'b000000000000000000110101000000
                ;mem[4681] <= 30'b000000000000000000110101010000
                ;mem[4682] <= 30'b000000000000000000110101100000
                ;mem[4683] <= 30'b000000000000000000110101110000
                ;mem[4684] <= 30'b000000000000000000110110000000
                ;mem[4685] <= 30'b000000000000000000110110010000
                ;mem[4686] <= 30'b000000000000000000111010010000
                ;mem[4687] <= 30'b000000000000000000111010100000
                ;mem[4688] <= 30'b000000000000000000111010110000
                ;mem[4689] <= 30'b000000000000000000111011000000
                ;mem[4690] <= 30'b000000000000000000111011010000
                ;mem[4691] <= 30'b000000000000000000111011100000
                ;mem[4692] <= 30'b000000000000000000111011110000
                ;mem[4693] <= 30'b000000000000000000111100000000
                ;mem[4694] <= 30'b000000000000000000111100010000
                ;mem[4695] <= 30'b000000000000000000111100100000
                ;mem[4696] <= 30'b000000000000000000111100110000
                ;mem[4697] <= 30'b000000000000000000111101000000
                ;mem[4698] <= 30'b000000000000000000111101010000
                ;mem[4699] <= 30'b000000001000000000000000000000
                ;mem[4700] <= 30'b000000001000000000000010110000
                ;mem[4701] <= 30'b000000001000000000000011000000
                ;mem[4702] <= 30'b000000001000000000000011010000
                ;mem[4703] <= 30'b000000001000000000000111000000
                ;mem[4704] <= 30'b000000001000000000000111010000
                ;mem[4705] <= 30'b000000001000000000000111100000
                ;mem[4706] <= 30'b000000001000000000000111110000
                ;mem[4707] <= 30'b000000001000000000001000000000
                ;mem[4708] <= 30'b000000001000000000001000010000
                ;mem[4709] <= 30'b000000001000000000001000100000
                ;mem[4710] <= 30'b000000001000000000001000110000
                ;mem[4711] <= 30'b000000001000000000001001000000
                ;mem[4712] <= 30'b000000001000000000001001010000
                ;mem[4713] <= 30'b000000001000000000001001100000
                ;mem[4714] <= 30'b000000001000000000001001110000
                ;mem[4715] <= 30'b000000001000000000001010000000
                ;mem[4716] <= 30'b000000001000000000001010010000
                ;mem[4717] <= 30'b000000001000000000001110010000
                ;mem[4718] <= 30'b000000001000000000001110100000
                ;mem[4719] <= 30'b000000001000000000001110110000
                ;mem[4720] <= 30'b000000001000000000001111000000
                ;mem[4721] <= 30'b000000001000000000001111010000
                ;mem[4722] <= 30'b000000001000000000001111100000
                ;mem[4723] <= 30'b000000001000000000001111110000
                ;mem[4724] <= 30'b000000001000000000010000000000
                ;mem[4725] <= 30'b000000001000000000010000010000
                ;mem[4726] <= 30'b000000001000000000010000100000
                ;mem[4727] <= 30'b000000001000000000010000110000
                ;mem[4728] <= 30'b000000001000000000010001000000
                ;mem[4729] <= 30'b000000001000000000010001010000
                ;mem[4730] <= 30'b000000001000000000010111100000
                ;mem[4731] <= 30'b000000001000000000010111110000
                ;mem[4732] <= 30'b000000001000000000011000000000
                ;mem[4733] <= 30'b000000001000000000011000010000
                ;mem[4734] <= 30'b000000001000000000011110100000
                ;mem[4735] <= 30'b000000001000000000011110110000
                ;mem[4736] <= 30'b000000001000000000011111000000
                ;mem[4737] <= 30'b000000001000000000100101100000
                ;mem[4738] <= 30'b000000001000000000100101110000
                ;mem[4739] <= 30'b000000001000000000100110000000
                ;mem[4740] <= 30'b000000001000000000101100010000
                ;mem[4741] <= 30'b000000001000000000101100100000
                ;mem[4742] <= 30'b000000001000000000101100110000
                ;mem[4743] <= 30'b000000001000000000101101000000
                ;mem[4744] <= 30'b000000001000000000110011000000
                ;mem[4745] <= 30'b000000001000000000110011010000
                ;mem[4746] <= 30'b000000001000000000110011100000
                ;mem[4747] <= 30'b000000001000000000111001110000
                ;mem[4748] <= 30'b000000001000000000111010000000
                ;mem[4749] <= 30'b000000001000000000111010010000
                ;mem[4750] <= 30'b000000001000000000111010100000
                ;mem[4751] <= 30'b000000010000000000000000010000
                ;mem[4752] <= 30'b000000010000000000000000100000
                ;mem[4753] <= 30'b000000010000000000000000110000
                ;mem[4754] <= 30'b000000010000000000000001000000
                ;mem[4755] <= 30'b000000010000000000000111000000
                ;mem[4756] <= 30'b000000010000000000000111010000
                ;mem[4757] <= 30'b000000010000000000000111100000
                ;mem[4758] <= 30'b000000010000000000001101110000
                ;mem[4759] <= 30'b000000010000000000001110000000
                ;mem[4760] <= 30'b000000010000000000001110010000
                ;mem[4761] <= 30'b000000010000000000001110100000
                ;mem[4762] <= 30'b000000010000000000010100100000
                ;mem[4763] <= 30'b000000010000000000010100110000
                ;mem[4764] <= 30'b000000010000000000010101000000
                ;mem[4765] <= 30'b000000010000000000010101010000
                ;mem[4766] <= 30'b000000010000000000011011010000
                ;mem[4767] <= 30'b000000010000000000011011100000
                ;mem[4768] <= 30'b000000010000000000011011110000
                ;mem[4769] <= 30'b000000010000000000011100000000
                ;mem[4770] <= 30'b000000010000000000011100010000
                ;mem[4771] <= 30'b000000010000000000100010010000
                ;mem[4772] <= 30'b000000010000000000100010100000
                ;mem[4773] <= 30'b000000010000000000100010110000
                ;mem[4774] <= 30'b000000010000000000100011000000
                ;mem[4775] <= 30'b000000010000000000101001000000
                ;mem[4776] <= 30'b000000010000000000101001010000
                ;mem[4777] <= 30'b000000010000000000101001100000
                ;mem[4778] <= 30'b000000010000000000101001110000
                ;mem[4779] <= 30'b000000010000000000101111110000
                ;mem[4780] <= 30'b000000010000000000110000000000
                ;mem[4781] <= 30'b000000010000000000110000010000
                ;mem[4782] <= 30'b000000010000000000110000100000
                ;mem[4783] <= 30'b000000010000000000110110100000
                ;mem[4784] <= 30'b000000010000000000110110110000
                ;mem[4785] <= 30'b000000010000000000110111000000
                ;mem[4786] <= 30'b000000010000000000110111010000
                ;mem[4787] <= 30'b000000010000000000111101100000
                ;mem[4788] <= 30'b000000010000000000111101110000
                ;mem[4789] <= 30'b000000010000000000111110000000
                ;mem[4790] <= 30'b000000010000000000111110010000
                ;mem[4791] <= 30'b000000000000000001000011110000
                ;mem[4792] <= 30'b000000000000000001000100000000
                ;mem[4793] <= 30'b000000000000000001000100010000
                ;mem[4794] <= 30'b000000000000000001000100100000
                ;mem[4795] <= 30'b000000000000000001001010100000
                ;mem[4796] <= 30'b000000000000000001001010110000
                ;mem[4797] <= 30'b000000000000000001001011000000
                ;mem[4798] <= 30'b000000000000000001001011010000
                ;mem[4799] <= 30'b000000000000000001010001100000
                ;mem[4800] <= 30'b000000000000000001010001110000
                ;mem[4801] <= 30'b000000000000000001010010000000
                ;mem[4802] <= 30'b000000000000000001010010010000
                ;mem[4803] <= 30'b000000000000000001011000000000
                ;mem[4804] <= 30'b000000000000000001011000010000
                ;mem[4805] <= 30'b000000000000000001011000100000
                ;mem[4806] <= 30'b000000000000000001011000110000
                ;mem[4807] <= 30'b000000000000000001011001000000
                ;mem[4808] <= 30'b000000000000000001011111000000
                ;mem[4809] <= 30'b000000000000000001011111010000
                ;mem[4810] <= 30'b000000000000000001011111100000
                ;mem[4811] <= 30'b000000000000000001011111110000
                ;mem[4812] <= 30'b000000000000000001100000000000
                ;mem[4813] <= 30'b000000000000000001100110000000
                ;mem[4814] <= 30'b000000000000000001100110010000
                ;mem[4815] <= 30'b000000000000000001100110100000
                ;mem[4816] <= 30'b000000000000000001100110110000
                ;mem[4817] <= 30'b000000000000000001101101000000
                ;mem[4818] <= 30'b000000000000000001101101010000
                ;mem[4819] <= 30'b000000000000000001101101100000
                ;mem[4820] <= 30'b000000000000000000011111100000
                ;mem[4821] <= 30'b000000000000000000011111110000
                ;mem[4822] <= 30'b000000000000000000100000000000
                ;mem[4823] <= 30'b000000000000000000100000010000
                ;mem[4824] <= 30'b000000000000000000100000100000
                ;mem[4825] <= 30'b000000000000000000100000110000
                ;mem[4826] <= 30'b000000000000000000100101110000
                ;mem[4827] <= 30'b000000000000000000100110000000
                ;mem[4828] <= 30'b000000000000000000100110010000
                ;mem[4829] <= 30'b000000000000000000100110100000
                ;mem[4830] <= 30'b000000000000000000100110110000
                ;mem[4831] <= 30'b000000000000000000100111000000
                ;mem[4832] <= 30'b000000000000000000100111010000
                ;mem[4833] <= 30'b000000000000000000100111100000
                ;mem[4834] <= 30'b000000000000000000100111110000
                ;mem[4835] <= 30'b000000000000000000101000000000
                ;mem[4836] <= 30'b000000000000000000101000010000
                ;mem[4837] <= 30'b000000000000000000101100100000
                ;mem[4838] <= 30'b000000000000000000101100110000
                ;mem[4839] <= 30'b000000000000000000101101000000
                ;mem[4840] <= 30'b000000000000000000101101010000
                ;mem[4841] <= 30'b000000000000000000101101100000
                ;mem[4842] <= 30'b000000000000000000101111000000
                ;mem[4843] <= 30'b000000000000000000101111010000
                ;mem[4844] <= 30'b000000000000000000110011010000
                ;mem[4845] <= 30'b000000000000000000110011100000
                ;mem[4846] <= 30'b000000000000000000110011110000
                ;mem[4847] <= 30'b000000000000000000110110000000
                ;mem[4848] <= 30'b000000000000000000110110010000
                ;mem[4849] <= 30'b000000000000000000111010000000
                ;mem[4850] <= 30'b000000000000000000111010010000
                ;mem[4851] <= 30'b000000000000000000111010100000
                ;mem[4852] <= 30'b000000000000000000111101000000
                ;mem[4853] <= 30'b000000000000000000111101010000
                ;mem[4854] <= 30'b000000001000000000000000100000
                ;mem[4855] <= 30'b000000001000000000000000110000
                ;mem[4856] <= 30'b000000001000000000000001000000
                ;mem[4857] <= 30'b000000001000000000000001010000
                ;mem[4858] <= 30'b000000001000000000000001100000
                ;mem[4859] <= 30'b000000001000000000000011000000
                ;mem[4860] <= 30'b000000001000000000000011010000
                ;mem[4861] <= 30'b000000001000000000000111010000
                ;mem[4862] <= 30'b000000001000000000000111100000
                ;mem[4863] <= 30'b000000001000000000000111110000
                ;mem[4864] <= 30'b000000001000000000001010000000
                ;mem[4865] <= 30'b000000001000000000001010010000
                ;mem[4866] <= 30'b000000001000000000001110000000
                ;mem[4867] <= 30'b000000001000000000001110010000
                ;mem[4868] <= 30'b000000001000000000001110100000
                ;mem[4869] <= 30'b000000001000000000010001000000
                ;mem[4870] <= 30'b000000001000000000010001010000
                ;mem[4871] <= 30'b000000001000000000010100110000
                ;mem[4872] <= 30'b000000001000000000010101000000
                ;mem[4873] <= 30'b000000001000000000011000000000
                ;mem[4874] <= 30'b000000001000000000011000010000
                ;mem[4875] <= 30'b000000001000000000011011110000
                ;mem[4876] <= 30'b000000001000000000011111000000
                ;mem[4877] <= 30'b000000001000000000011111010000
                ;mem[4878] <= 30'b000000001000000000100110000000
                ;mem[4879] <= 30'b000000001000000000100110010000
                ;mem[4880] <= 30'b000000001000000000101100110000
                ;mem[4881] <= 30'b000000001000000000101101000000
                ;mem[4882] <= 30'b000000001000000000110011100000
                ;mem[4883] <= 30'b000000001000000000110011110000
                ;mem[4884] <= 30'b000000001000000000110100000000
                ;mem[4885] <= 30'b000000001000000000111010010000
                ;mem[4886] <= 30'b000000001000000000111010100000
                ;mem[4887] <= 30'b000000001000000000111010110000
                ;mem[4888] <= 30'b000000010000000000000000110000
                ;mem[4889] <= 30'b000000010000000000000001000000
                ;mem[4890] <= 30'b000000010000000000000111100000
                ;mem[4891] <= 30'b000000010000000000000111110000
                ;mem[4892] <= 30'b000000010000000000001000000000
                ;mem[4893] <= 30'b000000010000000000001110010000
                ;mem[4894] <= 30'b000000010000000000001110100000
                ;mem[4895] <= 30'b000000010000000000001110110000
                ;mem[4896] <= 30'b000000010000000000010101000000
                ;mem[4897] <= 30'b000000010000000000010101010000
                ;mem[4898] <= 30'b000000010000000000010101100000
                ;mem[4899] <= 30'b000000010000000000011011110000
                ;mem[4900] <= 30'b000000010000000000011100000000
                ;mem[4901] <= 30'b000000010000000000011100010000
                ;mem[4902] <= 30'b000000010000000000100010100000
                ;mem[4903] <= 30'b000000010000000000100010110000
                ;mem[4904] <= 30'b000000010000000000100011000000
                ;mem[4905] <= 30'b000000010000000000101000110000
                ;mem[4906] <= 30'b000000010000000000101001000000
                ;mem[4907] <= 30'b000000010000000000101001010000
                ;mem[4908] <= 30'b000000010000000000101001100000
                ;mem[4909] <= 30'b000000010000000000101001110000
                ;mem[4910] <= 30'b000000010000000000101111000000
                ;mem[4911] <= 30'b000000010000000000101111010000
                ;mem[4912] <= 30'b000000010000000000101111100000
                ;mem[4913] <= 30'b000000010000000000101111110000
                ;mem[4914] <= 30'b000000010000000000110000000000
                ;mem[4915] <= 30'b000000010000000000110000010000
                ;mem[4916] <= 30'b000000010000000000110000100000
                ;mem[4917] <= 30'b000000010000000000110000110000
                ;mem[4918] <= 30'b000000010000000000110001000000
                ;mem[4919] <= 30'b000000010000000000110010100000
                ;mem[4920] <= 30'b000000010000000000110101100000
                ;mem[4921] <= 30'b000000010000000000110101110000
                ;mem[4922] <= 30'b000000010000000000110110000000
                ;mem[4923] <= 30'b000000010000000000110110010000
                ;mem[4924] <= 30'b000000010000000000110110100000
                ;mem[4925] <= 30'b000000010000000000110110110000
                ;mem[4926] <= 30'b000000010000000000110111000000
                ;mem[4927] <= 30'b000000010000000000110111010000
                ;mem[4928] <= 30'b000000010000000000110111100000
                ;mem[4929] <= 30'b000000010000000000110111110000
                ;mem[4930] <= 30'b000000010000000000111000000000
                ;mem[4931] <= 30'b000000010000000000111000010000
                ;mem[4932] <= 30'b000000010000000000111000100000
                ;mem[4933] <= 30'b000000010000000000111000110000
                ;mem[4934] <= 30'b000000010000000000111001010000
                ;mem[4935] <= 30'b000000010000000000111100010000
                ;mem[4936] <= 30'b000000010000000000111100100000
                ;mem[4937] <= 30'b000000010000000000111100110000
                ;mem[4938] <= 30'b000000010000000000111101000000
                ;mem[4939] <= 30'b000000010000000000111101010000
                ;mem[4940] <= 30'b000000010000000000111101100000
                ;mem[4941] <= 30'b000000010000000000111101110000
                ;mem[4942] <= 30'b000000010000000000111111000000
                ;mem[4943] <= 30'b000000010000000000111111010000
                ;mem[4944] <= 30'b000000010000000000111111100000
                ;mem[4945] <= 30'b000000010000000000111111110000
                ;mem[4946] <= 30'b000000000000000001000011000000
                ;mem[4947] <= 30'b000000000000000001000011010000
                ;mem[4948] <= 30'b000000000000000001000011100000
                ;mem[4949] <= 30'b000000000000000001000011110000
                ;mem[4950] <= 30'b000000000000000001000100000000
                ;mem[4951] <= 30'b000000000000000001000100010000
                ;mem[4952] <= 30'b000000000000000001000100100000
                ;mem[4953] <= 30'b000000000000000001000100110000
                ;mem[4954] <= 30'b000000000000000001000101000000
                ;mem[4955] <= 30'b000000000000000001000110100000
                ;mem[4956] <= 30'b000000000000000001001001100000
                ;mem[4957] <= 30'b000000000000000001001001110000
                ;mem[4958] <= 30'b000000000000000001001010000000
                ;mem[4959] <= 30'b000000000000000001001010010000
                ;mem[4960] <= 30'b000000000000000001001010100000
                ;mem[4961] <= 30'b000000000000000001001010110000
                ;mem[4962] <= 30'b000000000000000001001011000000
                ;mem[4963] <= 30'b000000000000000001001011010000
                ;mem[4964] <= 30'b000000000000000001001011100000
                ;mem[4965] <= 30'b000000000000000001001011110000
                ;mem[4966] <= 30'b000000000000000001001100000000
                ;mem[4967] <= 30'b000000000000000001001100010000
                ;mem[4968] <= 30'b000000000000000001001100100000
                ;mem[4969] <= 30'b000000000000000001001100110000
                ;mem[4970] <= 30'b000000000000000001001101010000
                ;mem[4971] <= 30'b000000000000000001010000010000
                ;mem[4972] <= 30'b000000000000000001010000100000
                ;mem[4973] <= 30'b000000000000000001010000110000
                ;mem[4974] <= 30'b000000000000000001010001000000
                ;mem[4975] <= 30'b000000000000000001010001010000
                ;mem[4976] <= 30'b000000000000000001010001100000
                ;mem[4977] <= 30'b000000000000000001010001110000
                ;mem[4978] <= 30'b000000000000000001010011000000
                ;mem[4979] <= 30'b000000000000000001010011010000
                ;mem[4980] <= 30'b000000000000000001010011100000
                ;mem[4981] <= 30'b000000000000000001010011110000
                ;mem[4982] <= 30'b000000000000000001010100000000
                ;mem[4983] <= 30'b000000000000000001010100010000
                ;mem[4984] <= 30'b000000000000000001010111010000
                ;mem[4985] <= 30'b000000000000000001010111100000
                ;mem[4986] <= 30'b000000000000000001010111110000
                ;mem[4987] <= 30'b000000000000000001011000000000
                ;mem[4988] <= 30'b000000000000000001011000010000
                ;mem[4989] <= 30'b000000000000000001011000100000
                ;mem[4990] <= 30'b000000000000000001011010100000
                ;mem[4991] <= 30'b000000000000000001011010110000
                ;mem[4992] <= 30'b000000000000000001011110110000
                ;mem[4993] <= 30'b000000000000000001011111000000
                ;mem[4994] <= 30'b000000000000000000110010110000
                ;mem[4995] <= 30'b000000000000000000110011000000
                ;mem[4996] <= 30'b000000000000000000110011110000
                ;mem[4997] <= 30'b000000000000000000110100000000
                ;mem[4998] <= 30'b000000000000000000110100010000
                ;mem[4999] <= 30'b000000000000000000110100100000
                ;mem[5000] <= 30'b000000000000000000110100110000
                ;mem[5001] <= 30'b000000000000000000110101000000
                ;mem[5002] <= 30'b000000000000000000110101010000
                ;mem[5003] <= 30'b000000000000000000110101100000
                ;mem[5004] <= 30'b000000000000000000111001100000
                ;mem[5005] <= 30'b000000000000000000111001110000
                ;mem[5006] <= 30'b000000000000000000111010000000
                ;mem[5007] <= 30'b000000000000000000111010010000
                ;mem[5008] <= 30'b000000000000000000111010100000
                ;mem[5009] <= 30'b000000000000000000111010110000
                ;mem[5010] <= 30'b000000000000000000111011000000
                ;mem[5011] <= 30'b000000000000000000111011010000
                ;mem[5012] <= 30'b000000000000000000111011100000
                ;mem[5013] <= 30'b000000000000000000111011110000
                ;mem[5014] <= 30'b000000000000000000111100000000
                ;mem[5015] <= 30'b000000000000000000111100010000
                ;mem[5016] <= 30'b000000000000000000111100100000
                ;mem[5017] <= 30'b000000000000000000111100110000
                ;mem[5018] <= 30'b000000001000000000000110110000
                ;mem[5019] <= 30'b000000001000000000000111000000
                ;mem[5020] <= 30'b000000001000000000000111110000
                ;mem[5021] <= 30'b000000001000000000001000000000
                ;mem[5022] <= 30'b000000001000000000001000010000
                ;mem[5023] <= 30'b000000001000000000001000100000
                ;mem[5024] <= 30'b000000001000000000001000110000
                ;mem[5025] <= 30'b000000001000000000001001000000
                ;mem[5026] <= 30'b000000001000000000001001010000
                ;mem[5027] <= 30'b000000001000000000001001100000
                ;mem[5028] <= 30'b000000001000000000001101100000
                ;mem[5029] <= 30'b000000001000000000001101110000
                ;mem[5030] <= 30'b000000001000000000001110000000
                ;mem[5031] <= 30'b000000001000000000001110010000
                ;mem[5032] <= 30'b000000001000000000001110100000
                ;mem[5033] <= 30'b000000001000000000001110110000
                ;mem[5034] <= 30'b000000001000000000001111000000
                ;mem[5035] <= 30'b000000001000000000001111010000
                ;mem[5036] <= 30'b000000001000000000001111100000
                ;mem[5037] <= 30'b000000001000000000001111110000
                ;mem[5038] <= 30'b000000001000000000010000000000
                ;mem[5039] <= 30'b000000001000000000010000010000
                ;mem[5040] <= 30'b000000001000000000010000100000
                ;mem[5041] <= 30'b000000001000000000010000110000
                ;mem[5042] <= 30'b000000001000000000010100010000
                ;mem[5043] <= 30'b000000001000000000010100100000
                ;mem[5044] <= 30'b000000001000000000010100110000
                ;mem[5045] <= 30'b000000001000000000010101000000
                ;mem[5046] <= 30'b000000001000000000010101010000
                ;mem[5047] <= 30'b000000001000000000010101100000
                ;mem[5048] <= 30'b000000001000000000010111100000
                ;mem[5049] <= 30'b000000001000000000010111110000
                ;mem[5050] <= 30'b000000001000000000011011000000
                ;mem[5051] <= 30'b000000001000000000011011010000
                ;mem[5052] <= 30'b000000001000000000011011100000
                ;mem[5053] <= 30'b000000001000000000011011110000
                ;mem[5054] <= 30'b000000001000000000011110100000
                ;mem[5055] <= 30'b000000001000000000011110110000
                ;mem[5056] <= 30'b000000001000000000100001110000
                ;mem[5057] <= 30'b000000001000000000100010000000
                ;mem[5058] <= 30'b000000001000000000100010010000
                ;mem[5059] <= 30'b000000001000000000100010100000
                ;mem[5060] <= 30'b000000001000000000100101100000
                ;mem[5061] <= 30'b000000001000000000100101110000
                ;mem[5062] <= 30'b000000001000000000101000110000
                ;mem[5063] <= 30'b000000001000000000101001000000
                ;mem[5064] <= 30'b000000001000000000101100010000
                ;mem[5065] <= 30'b000000001000000000101100100000
                ;mem[5066] <= 30'b000000001000000000101100110000
                ;mem[5067] <= 30'b000000001000000000110011010000
                ;mem[5068] <= 30'b000000001000000000110011100000
                ;mem[5069] <= 30'b000000001000000000111010000000
                ;mem[5070] <= 30'b000000001000000000111010010000
                ;mem[5071] <= 30'b000000001000000000111010100000
                ;mem[5072] <= 30'b000000010000000000000000010000
                ;mem[5073] <= 30'b000000010000000000000000100000
                ;mem[5074] <= 30'b000000010000000000000000110000
                ;mem[5075] <= 30'b000000010000000000000111010000
                ;mem[5076] <= 30'b000000010000000000000111100000
                ;mem[5077] <= 30'b000000010000000000001110000000
                ;mem[5078] <= 30'b000000010000000000001110010000
                ;mem[5079] <= 30'b000000010000000000001110100000
                ;mem[5080] <= 30'b000000010000000000010101000000
                ;mem[5081] <= 30'b000000010000000000010101010000
                ;mem[5082] <= 30'b000000010000000000011100000000
                ;mem[5083] <= 30'b000000010000000000011100010000
                ;mem[5084] <= 30'b000000010000000000100010110000
                ;mem[5085] <= 30'b000000010000000000100011000000
                ;mem[5086] <= 30'b000000010000000000101001110000
                ;mem[5087] <= 30'b000000010000000000101010000000
                ;mem[5088] <= 30'b000000010000000000101010010000
                ;mem[5089] <= 30'b000000010000000000101010100000
                ;mem[5090] <= 30'b000000010000000000101010110000
                ;mem[5091] <= 30'b000000010000000000101011000000
                ;mem[5092] <= 30'b000000010000000000110000010000
                ;mem[5093] <= 30'b000000010000000000110000100000
                ;mem[5094] <= 30'b000000010000000000110000110000
                ;mem[5095] <= 30'b000000010000000000110001000000
                ;mem[5096] <= 30'b000000010000000000110001010000
                ;mem[5097] <= 30'b000000010000000000110001100000
                ;mem[5098] <= 30'b000000010000000000110001110000
                ;mem[5099] <= 30'b000000010000000000110010000000
                ;mem[5100] <= 30'b000000010000000000110111000000
                ;mem[5101] <= 30'b000000010000000000110111010000
                ;mem[5102] <= 30'b000000010000000000110111100000
                ;mem[5103] <= 30'b000000010000000000110111110000
                ;mem[5104] <= 30'b000000010000000000111000000000
                ;mem[5105] <= 30'b000000010000000000111110100000
                ;mem[5106] <= 30'b000000010000000000111110110000
                ;mem[5107] <= 30'b000000000000000001000100010000
                ;mem[5108] <= 30'b000000000000000001000100100000
                ;mem[5109] <= 30'b000000000000000001000100110000
                ;mem[5110] <= 30'b000000000000000001000101000000
                ;mem[5111] <= 30'b000000000000000001000101010000
                ;mem[5112] <= 30'b000000000000000001000101100000
                ;mem[5113] <= 30'b000000000000000001000101110000
                ;mem[5114] <= 30'b000000000000000001000110000000
                ;mem[5115] <= 30'b000000000000000001001011000000
                ;mem[5116] <= 30'b000000000000000001001011010000
                ;mem[5117] <= 30'b000000000000000001001011100000
                ;mem[5118] <= 30'b000000000000000001001011110000
                ;mem[5119] <= 30'b000000000000000001001100000000
                ;mem[5120] <= 30'b000000000000000001010010100000
                ;mem[5121] <= 30'b000000000000000001010010110000
                ;mem[5122] <= 30'b000000000000000001011001100000
                ;mem[5123] <= 30'b000000000000000001011001110000
                ;mem[5124] <= 30'b000000000000000001100000100000
                ;mem[5125] <= 30'b000000000000000001100000110000
                ;mem[5126] <= 30'b000000000000000001100111100000
                ;mem[5127] <= 30'b000000000000000001101110100000
                ;mem[5128] <= 30'b000000000000000001110101100000
                ;mem[5129] <= 30'b000000000000000000100110000000
                ;mem[5130] <= 30'b000000000000000000100110010000
                ;mem[5131] <= 30'b000000000000000000101101000000
                ;mem[5132] <= 30'b000000000000000000101101010000
                ;mem[5133] <= 30'b000000000000000000101101100000
                ;mem[5134] <= 30'b000000000000000000110100000000
                ;mem[5135] <= 30'b000000000000000000110100010000
                ;mem[5136] <= 30'b000000000000000000110100100000
                ;mem[5137] <= 30'b000000000000000000111011000000
                ;mem[5138] <= 30'b000000000000000000111011010000
                ;mem[5139] <= 30'b000000000000000000111011100000
                ;mem[5140] <= 30'b000000001000000000000001000000
                ;mem[5141] <= 30'b000000001000000000000001010000
                ;mem[5142] <= 30'b000000001000000000000001100000
                ;mem[5143] <= 30'b000000001000000000001000000000
                ;mem[5144] <= 30'b000000001000000000001000010000
                ;mem[5145] <= 30'b000000001000000000001000100000
                ;mem[5146] <= 30'b000000001000000000001111000000
                ;mem[5147] <= 30'b000000001000000000001111010000
                ;mem[5148] <= 30'b000000001000000000001111100000
                ;mem[5149] <= 30'b000000001000000000010110000000
                ;mem[5150] <= 30'b000000001000000000010110010000
                ;mem[5151] <= 30'b000000001000000000010110100000
                ;mem[5152] <= 30'b000000001000000000011101010000
                ;mem[5153] <= 30'b000000001000000000011101100000
                ;mem[5154] <= 30'b000000001000000000011101110000
                ;mem[5155] <= 30'b000000001000000000100100010000
                ;mem[5156] <= 30'b000000001000000000100100100000
                ;mem[5157] <= 30'b000000001000000000100100110000
                ;mem[5158] <= 30'b000000001000000000101011010000
                ;mem[5159] <= 30'b000000001000000000101011100000
                ;mem[5160] <= 30'b000000001000000000101011110000
                ;mem[5161] <= 30'b000000001000000000110010010000
                ;mem[5162] <= 30'b000000001000000000110010100000
                ;mem[5163] <= 30'b000000001000000000110010110000
                ;mem[5164] <= 30'b000000001000000000111001010000
                ;mem[5165] <= 30'b000000001000000000111001100000
                ;mem[5166] <= 30'b000000001000000000111001110000
                ;mem[5167] <= 30'b000000010000000000000110010000
                ;mem[5168] <= 30'b000000010000000000000110100000
                ;mem[5169] <= 30'b000000010000000000000110110000
                ;mem[5170] <= 30'b000000010000000000001101010000
                ;mem[5171] <= 30'b000000010000000000001101100000
                ;mem[5172] <= 30'b000000010000000000001101110000
                ;mem[5173] <= 30'b000000010000000000010100010000
                ;mem[5174] <= 30'b000000010000000000010100100000
                ;mem[5175] <= 30'b000000010000000000010100110000
                ;mem[5176] <= 30'b000000010000000000011011010000
                ;mem[5177] <= 30'b000000010000000000011011100000
                ;mem[5178] <= 30'b000000010000000000011011110000
                ;mem[5179] <= 30'b000000010000000000100010010000
                ;mem[5180] <= 30'b000000010000000000100010100000
                ;mem[5181] <= 30'b000000010000000000100010110000
                ;mem[5182] <= 30'b000000010000000000101001010000
                ;mem[5183] <= 30'b000000010000000000101001100000
                ;mem[5184] <= 30'b000000010000000000101001110000
                ;mem[5185] <= 30'b000000010000000000110000010000
                ;mem[5186] <= 30'b000000010000000000110000100000
                ;mem[5187] <= 30'b000000010000000000110000110000
                ;mem[5188] <= 30'b000000010000000000110111010000
                ;mem[5189] <= 30'b000000010000000000110111100000
                ;mem[5190] <= 30'b000000010000000000110111110000
                ;mem[5191] <= 30'b000000010000000000111110010000
                ;mem[5192] <= 30'b000000010000000000111110100000
                ;mem[5193] <= 30'b000000010000000000111110110000
                ;mem[5194] <= 30'b000000000000000001000100010000
                ;mem[5195] <= 30'b000000000000000001000100100000
                ;mem[5196] <= 30'b000000000000000001000100110000
                ;mem[5197] <= 30'b000000000000000001001011010000
                ;mem[5198] <= 30'b000000000000000001001011100000
                ;mem[5199] <= 30'b000000000000000001001011110000
                ;mem[5200] <= 30'b000000000000000001010010010000
                ;mem[5201] <= 30'b000000000000000001010010100000
                ;mem[5202] <= 30'b000000000000000001010010110000
                ;mem[5203] <= 30'b000000000000000001011001100000
                ;mem[5204] <= 30'b000000000000000001011001110000
                ;mem[5205] <= 30'b000000000000000001100000100000
                ;mem[5206] <= 30'b000000000000000001100000110000
                ;mem[5207] <= 30'b000000000000000001100111100000
                ;mem[5208] <= 30'b000000000000000001100111110000
                ;mem[5209] <= 30'b000000000000000000011111100000
                ;mem[5210] <= 30'b000000000000000000011111110000
                ;mem[5211] <= 30'b000000000000000000100110000000
                ;mem[5212] <= 30'b000000000000000000100110010000
                ;mem[5213] <= 30'b000000000000000000100110100000
                ;mem[5214] <= 30'b000000000000000000100110110000
                ;mem[5215] <= 30'b000000000000000000100111000000
                ;mem[5216] <= 30'b000000000000000000101100110000
                ;mem[5217] <= 30'b000000000000000000101101000000
                ;mem[5218] <= 30'b000000000000000000101101010000
                ;mem[5219] <= 30'b000000000000000000101101100000
                ;mem[5220] <= 30'b000000000000000000101101110000
                ;mem[5221] <= 30'b000000000000000000101110000000
                ;mem[5222] <= 30'b000000000000000000110011010000
                ;mem[5223] <= 30'b000000000000000000110011100000
                ;mem[5224] <= 30'b000000000000000000110011110000
                ;mem[5225] <= 30'b000000000000000000110100110000
                ;mem[5226] <= 30'b000000000000000000110101000000
                ;mem[5227] <= 30'b000000000000000000111010000000
                ;mem[5228] <= 30'b000000000000000000111010010000
                ;mem[5229] <= 30'b000000000000000000111011110000
                ;mem[5230] <= 30'b000000000000000000111100000000
                ;mem[5231] <= 30'b000000001000000000000000110000
                ;mem[5232] <= 30'b000000001000000000000001000000
                ;mem[5233] <= 30'b000000001000000000000001010000
                ;mem[5234] <= 30'b000000001000000000000001100000
                ;mem[5235] <= 30'b000000001000000000000001110000
                ;mem[5236] <= 30'b000000001000000000000010000000
                ;mem[5237] <= 30'b000000001000000000000111010000
                ;mem[5238] <= 30'b000000001000000000000111100000
                ;mem[5239] <= 30'b000000001000000000000111110000
                ;mem[5240] <= 30'b000000001000000000001000110000
                ;mem[5241] <= 30'b000000001000000000001001000000
                ;mem[5242] <= 30'b000000001000000000001110000000
                ;mem[5243] <= 30'b000000001000000000001110010000
                ;mem[5244] <= 30'b000000001000000000001111110000
                ;mem[5245] <= 30'b000000001000000000010000000000
                ;mem[5246] <= 30'b000000001000000000010110110000
                ;mem[5247] <= 30'b000000001000000000011101110000
                ;mem[5248] <= 30'b000000001000000000100100100000
                ;mem[5249] <= 30'b000000001000000000100100110000
                ;mem[5250] <= 30'b000000001000000000101011010000
                ;mem[5251] <= 30'b000000001000000000101011100000
                ;mem[5252] <= 30'b000000001000000000110010010000
                ;mem[5253] <= 30'b000000001000000000110010100000
                ;mem[5254] <= 30'b000000001000000000111001000000
                ;mem[5255] <= 30'b000000001000000000111001010000
                ;mem[5256] <= 30'b000000010000000000000110010000
                ;mem[5257] <= 30'b000000010000000000000110100000
                ;mem[5258] <= 30'b000000010000000000001101000000
                ;mem[5259] <= 30'b000000010000000000001101010000
                ;mem[5260] <= 30'b000000010000000000010100000000
                ;mem[5261] <= 30'b000000010000000000010100010000
                ;mem[5262] <= 30'b000000010000000000011010110000
                ;mem[5263] <= 30'b000000010000000000011011000000
                ;mem[5264] <= 30'b000000010000000000011101110000
                ;mem[5265] <= 30'b000000010000000000100001110000
                ;mem[5266] <= 30'b000000010000000000100010000000
                ;mem[5267] <= 30'b000000010000000000100100010000
                ;mem[5268] <= 30'b000000010000000000100100100000
                ;mem[5269] <= 30'b000000010000000000100100110000
                ;mem[5270] <= 30'b000000010000000000101000100000
                ;mem[5271] <= 30'b000000010000000000101000110000
                ;mem[5272] <= 30'b000000010000000000101010100000
                ;mem[5273] <= 30'b000000010000000000101010110000
                ;mem[5274] <= 30'b000000010000000000101011000000
                ;mem[5275] <= 30'b000000010000000000101011010000
                ;mem[5276] <= 30'b000000010000000000101111010000
                ;mem[5277] <= 30'b000000010000000000101111100000
                ;mem[5278] <= 30'b000000010000000000110001000000
                ;mem[5279] <= 30'b000000010000000000110001010000
                ;mem[5280] <= 30'b000000010000000000110001100000
                ;mem[5281] <= 30'b000000010000000000110001110000
                ;mem[5282] <= 30'b000000010000000000110110010000
                ;mem[5283] <= 30'b000000010000000000110110100000
                ;mem[5284] <= 30'b000000010000000000110111100000
                ;mem[5285] <= 30'b000000010000000000110111110000
                ;mem[5286] <= 30'b000000010000000000111000000000
                ;mem[5287] <= 30'b000000010000000000111000010000
                ;mem[5288] <= 30'b000000010000000000111101000000
                ;mem[5289] <= 30'b000000010000000000111101010000
                ;mem[5290] <= 30'b000000010000000000111101110000
                ;mem[5291] <= 30'b000000010000000000111110000000
                ;mem[5292] <= 30'b000000010000000000111110010000
                ;mem[5293] <= 30'b000000010000000000111110100000
                ;mem[5294] <= 30'b000000010000000000111110110000
                ;mem[5295] <= 30'b000000000000000001000011010000
                ;mem[5296] <= 30'b000000000000000001000011100000
                ;mem[5297] <= 30'b000000000000000001000101000000
                ;mem[5298] <= 30'b000000000000000001000101010000
                ;mem[5299] <= 30'b000000000000000001000101100000
                ;mem[5300] <= 30'b000000000000000001000101110000
                ;mem[5301] <= 30'b000000000000000001001010010000
                ;mem[5302] <= 30'b000000000000000001001010100000
                ;mem[5303] <= 30'b000000000000000001001011100000
                ;mem[5304] <= 30'b000000000000000001001011110000
                ;mem[5305] <= 30'b000000000000000001001100000000
                ;mem[5306] <= 30'b000000000000000001001100010000
                ;mem[5307] <= 30'b000000000000000001010001000000
                ;mem[5308] <= 30'b000000000000000001010001010000
                ;mem[5309] <= 30'b000000000000000001010001110000
                ;mem[5310] <= 30'b000000000000000001010010000000
                ;mem[5311] <= 30'b000000000000000001010010010000
                ;mem[5312] <= 30'b000000000000000001010010100000
                ;mem[5313] <= 30'b000000000000000001010010110000
                ;mem[5314] <= 30'b000000000000000001011000000000
                ;mem[5315] <= 30'b000000000000000001011000010000
                ;mem[5316] <= 30'b000000000000000001011000100000
                ;mem[5317] <= 30'b000000000000000001011000110000
                ;mem[5318] <= 30'b000000000000000001011001000000
                ;mem[5319] <= 30'b000000000000000001011001010000
                ;mem[5320] <= 30'b000000000000000001011111000000
                ;mem[5321] <= 30'b000000000000000001011111010000
                ;mem[5322] <= 30'b000000000000000001011111100000
                ;mem[5323] <= 30'b000000000000000000011111110000
                ;mem[5324] <= 30'b000000000000000000100110100000
                ;mem[5325] <= 30'b000000000000000000100110110000
                ;mem[5326] <= 30'b000000000000000000101101100000
                ;mem[5327] <= 30'b000000000000000000101101110000
                ;mem[5328] <= 30'b000000000000000000101110000000
                ;mem[5329] <= 30'b000000000000000000101110010000
                ;mem[5330] <= 30'b000000000000000000110100010000
                ;mem[5331] <= 30'b000000000000000000110100100000
                ;mem[5332] <= 30'b000000000000000000110100110000
                ;mem[5333] <= 30'b000000000000000000110101000000
                ;mem[5334] <= 30'b000000000000000000110101010000
                ;mem[5335] <= 30'b000000000000000000111011010000
                ;mem[5336] <= 30'b000000000000000000111011100000
                ;mem[5337] <= 30'b000000000000000000111011110000
                ;mem[5338] <= 30'b000000000000000000111100000000
                ;mem[5339] <= 30'b000000000000000000111100010000
                ;mem[5340] <= 30'b000000001000000000000001100000
                ;mem[5341] <= 30'b000000001000000000000001110000
                ;mem[5342] <= 30'b000000001000000000000010000000
                ;mem[5343] <= 30'b000000001000000000000010010000
                ;mem[5344] <= 30'b000000001000000000001000010000
                ;mem[5345] <= 30'b000000001000000000001000100000
                ;mem[5346] <= 30'b000000001000000000001000110000
                ;mem[5347] <= 30'b000000001000000000001001000000
                ;mem[5348] <= 30'b000000001000000000001001010000
                ;mem[5349] <= 30'b000000001000000000001111010000
                ;mem[5350] <= 30'b000000001000000000001111100000
                ;mem[5351] <= 30'b000000001000000000001111110000
                ;mem[5352] <= 30'b000000001000000000010000000000
                ;mem[5353] <= 30'b000000001000000000010000010000
                ;mem[5354] <= 30'b000000001000000000010110010000
                ;mem[5355] <= 30'b000000001000000000010110100000
                ;mem[5356] <= 30'b000000001000000000010110110000
                ;mem[5357] <= 30'b000000001000000000010111000000
                ;mem[5358] <= 30'b000000001000000000011101010000
                ;mem[5359] <= 30'b000000001000000000011101100000
                ;mem[5360] <= 30'b000000001000000000011101110000
                ;mem[5361] <= 30'b000000001000000000011110000000
                ;mem[5362] <= 30'b000000001000000000100100000000
                ;mem[5363] <= 30'b000000001000000000100100010000
                ;mem[5364] <= 30'b000000001000000000100100100000
                ;mem[5365] <= 30'b000000001000000000100100110000
                ;mem[5366] <= 30'b000000001000000000100101000000
                ;mem[5367] <= 30'b000000001000000000101011000000
                ;mem[5368] <= 30'b000000001000000000101011010000
                ;mem[5369] <= 30'b000000001000000000101011100000
                ;mem[5370] <= 30'b000000001000000000101011110000
                ;mem[5371] <= 30'b000000001000000000110010000000
                ;mem[5372] <= 30'b000000001000000000110010010000
                ;mem[5373] <= 30'b000000001000000000110010100000
                ;mem[5374] <= 30'b000000001000000000110010110000
                ;mem[5375] <= 30'b000000001000000000111001000000
                ;mem[5376] <= 30'b000000001000000000111001010000
                ;mem[5377] <= 30'b000000001000000000111001100000
                ;mem[5378] <= 30'b000000001000000000111001110000
                ;mem[5379] <= 30'b000000010000000000000110000000
                ;mem[5380] <= 30'b000000010000000000000110010000
                ;mem[5381] <= 30'b000000010000000000000110100000
                ;mem[5382] <= 30'b000000010000000000000110110000
                ;mem[5383] <= 30'b000000010000000000001101000000
                ;mem[5384] <= 30'b000000010000000000001101010000
                ;mem[5385] <= 30'b000000010000000000001101100000
                ;mem[5386] <= 30'b000000010000000000001101110000
                ;mem[5387] <= 30'b000000010000000000010100000000
                ;mem[5388] <= 30'b000000010000000000010100010000
                ;mem[5389] <= 30'b000000010000000000010100100000
                ;mem[5390] <= 30'b000000010000000000010100110000
                ;mem[5391] <= 30'b000000010000000000011011000000
                ;mem[5392] <= 30'b000000010000000000011011010000
                ;mem[5393] <= 30'b000000010000000000011011100000
                ;mem[5394] <= 30'b000000010000000000100010000000
                ;mem[5395] <= 30'b000000010000000000100010010000
                ;mem[5396] <= 30'b000000010000000000100010100000
                ;mem[5397] <= 30'b000000010000000000101001000000
                ;mem[5398] <= 30'b000000010000000000101001010000
                ;mem[5399] <= 30'b000000010000000000101001100000
                ;mem[5400] <= 30'b000000010000000000110000000000
                ;mem[5401] <= 30'b000000010000000000110000010000
                ;mem[5402] <= 30'b000000010000000000110000100000
                ;mem[5403] <= 30'b000000010000000000110000110000
                ;mem[5404] <= 30'b000000010000000000110111000000
                ;mem[5405] <= 30'b000000010000000000110111010000
                ;mem[5406] <= 30'b000000010000000000110111100000
                ;mem[5407] <= 30'b000000010000000000110111110000
                ;mem[5408] <= 30'b000000010000000000111110000000
                ;mem[5409] <= 30'b000000010000000000111110010000
                ;mem[5410] <= 30'b000000010000000000111110100000
                ;mem[5411] <= 30'b000000010000000000111110110000
                ;mem[5412] <= 30'b000000000000000001000100000000
                ;mem[5413] <= 30'b000000000000000001000100010000
                ;mem[5414] <= 30'b000000000000000001000100100000
                ;mem[5415] <= 30'b000000000000000001000100110000
                ;mem[5416] <= 30'b000000000000000001001011000000
                ;mem[5417] <= 30'b000000000000000001001011010000
                ;mem[5418] <= 30'b000000000000000001001011100000
                ;mem[5419] <= 30'b000000000000000001001011110000
                ;mem[5420] <= 30'b000000000000000001010010000000
                ;mem[5421] <= 30'b000000000000000001010010010000
                ;mem[5422] <= 30'b000000000000000001010010100000
                ;mem[5423] <= 30'b000000000000000001010010110000
                ;mem[5424] <= 30'b000000000000000001011001000000
                ;mem[5425] <= 30'b000000000000000001011001010000
                ;mem[5426] <= 30'b000000000000000001011001100000
                ;mem[5427] <= 30'b000000000000000001011001110000
                ;mem[5428] <= 30'b000000000000000001100000010000
                ;mem[5429] <= 30'b000000000000000001100000100000
                ;mem[5430] <= 30'b000000000000000000011111010000
                ;mem[5431] <= 30'b000000000000000000100110010000
                ;mem[5432] <= 30'b000000000000000000100110100000
                ;mem[5433] <= 30'b000000000000000000101101010000
                ;mem[5434] <= 30'b000000000000000000101101100000
                ;mem[5435] <= 30'b000000000000000000110100100000
                ;mem[5436] <= 30'b000000000000000000111011100000
                ;mem[5437] <= 30'b000000001000000000000001010000
                ;mem[5438] <= 30'b000000001000000000000001100000
                ;mem[5439] <= 30'b000000001000000000001000100000
                ;mem[5440] <= 30'b000000001000000000001111100000
                ;mem[5441] <= 30'b000000001000000000010110100000
                ;mem[5442] <= 30'b000000001000000000011101100000
                ;mem[5443] <= 30'b000000001000000000100100100000
                ;mem[5444] <= 30'b000000001000000000101011100000
                ;mem[5445] <= 30'b000000001000000000110010100000
                ;mem[5446] <= 30'b000000001000000000111001100000
                ;mem[5447] <= 30'b000000010000000000000110100000
                ;mem[5448] <= 30'b000000010000000000001101100000
                ;mem[5449] <= 30'b000000010000000000010100100000
                ;mem[5450] <= 30'b000000010000000000011011100000
                ;mem[5451] <= 30'b000000010000000000100010010000
                ;mem[5452] <= 30'b000000010000000000100010100000
                ;mem[5453] <= 30'b000000010000000000101001010000
                ;mem[5454] <= 30'b000000010000000000101001100000
                ;mem[5455] <= 30'b000000010000000000110000010000
                ;mem[5456] <= 30'b000000010000000000110000100000
                ;mem[5457] <= 30'b000000010000000000110111010000
                ;mem[5458] <= 30'b000000010000000000110111100000
                ;mem[5459] <= 30'b000000010000000000111110010000
                ;mem[5460] <= 30'b000000000000000001000100010000
                ;mem[5461] <= 30'b000000000000000001000100100000
                ;mem[5462] <= 30'b000000000000000001001011010000
                ;mem[5463] <= 30'b000000000000000001001011100000
                ;mem[5464] <= 30'b000000000000000001010010010000
                ;mem[5465] <= 30'b000000000000000001011001010000
                ;mem[5466] <= 30'b000000000000000001100000010000
                ;mem[5467] <= 30'b000000000000000000110100010000
                ;mem[5468] <= 30'b000000000000000000110100100000
                ;mem[5469] <= 30'b000000000000000000110100110000
                ;mem[5470] <= 30'b000000000000000000110101000000
                ;mem[5471] <= 30'b000000000000000000111010010000
                ;mem[5472] <= 30'b000000000000000000111010100000
                ;mem[5473] <= 30'b000000000000000000111010110000
                ;mem[5474] <= 30'b000000000000000000111011000000
                ;mem[5475] <= 30'b000000000000000000111011010000
                ;mem[5476] <= 30'b000000000000000000111011100000
                ;mem[5477] <= 30'b000000000000000000111011110000
                ;mem[5478] <= 30'b000000000000000000111100000000
                ;mem[5479] <= 30'b000000000000000000111100010000
                ;mem[5480] <= 30'b000000001000000000001000010000
                ;mem[5481] <= 30'b000000001000000000001000100000
                ;mem[5482] <= 30'b000000001000000000001000110000
                ;mem[5483] <= 30'b000000001000000000001001000000
                ;mem[5484] <= 30'b000000001000000000001110010000
                ;mem[5485] <= 30'b000000001000000000001110100000
                ;mem[5486] <= 30'b000000001000000000001110110000
                ;mem[5487] <= 30'b000000001000000000001111000000
                ;mem[5488] <= 30'b000000001000000000001111010000
                ;mem[5489] <= 30'b000000001000000000001111100000
                ;mem[5490] <= 30'b000000001000000000001111110000
                ;mem[5491] <= 30'b000000001000000000010000000000
                ;mem[5492] <= 30'b000000001000000000010000010000
                ;mem[5493] <= 30'b000000001000000000010100110000
                ;mem[5494] <= 30'b000000001000000000010101000000
                ;mem[5495] <= 30'b000000001000000000010101010000
                ;mem[5496] <= 30'b000000001000000000010101100000
                ;mem[5497] <= 30'b000000001000000000010101110000
                ;mem[5498] <= 30'b000000001000000000010110000000
                ;mem[5499] <= 30'b000000001000000000010110010000
                ;mem[5500] <= 30'b000000001000000000010111000000
                ;mem[5501] <= 30'b000000001000000000010111010000
                ;mem[5502] <= 30'b000000001000000000011011110000
                ;mem[5503] <= 30'b000000001000000000011100000000
                ;mem[5504] <= 30'b000000001000000000011100010000
                ;mem[5505] <= 30'b000000001000000000011110010000
                ;mem[5506] <= 30'b000000001000000000100101010000
                ;mem[5507] <= 30'b000000001000000000100101100000
                ;mem[5508] <= 30'b000000001000000000101100010000
                ;mem[5509] <= 30'b000000001000000000101100100000
                ;mem[5510] <= 30'b000000001000000000110011010000
                ;mem[5511] <= 30'b000000001000000000111010000000
                ;mem[5512] <= 30'b000000001000000000111010010000
                ;mem[5513] <= 30'b000000010000000000000000010000
                ;mem[5514] <= 30'b000000010000000000000000100000
                ;mem[5515] <= 30'b000000010000000000000111010000
                ;mem[5516] <= 30'b000000010000000000001110000000
                ;mem[5517] <= 30'b000000010000000000001110010000
                ;mem[5518] <= 30'b000000010000000000010101000000
                ;mem[5519] <= 30'b000000010000000000011011100000
                ;mem[5520] <= 30'b000000010000000000011011110000
                ;mem[5521] <= 30'b000000010000000000011100000000
                ;mem[5522] <= 30'b000000010000000000100010100000
                ;mem[5523] <= 30'b000000010000000000100010110000
                ;mem[5524] <= 30'b000000010000000000100011000000
                ;mem[5525] <= 30'b000000010000000000100011010000
                ;mem[5526] <= 30'b000000010000000000100011100000
                ;mem[5527] <= 30'b000000010000000000100011110000
                ;mem[5528] <= 30'b000000010000000000101001100000
                ;mem[5529] <= 30'b000000010000000000101001110000
                ;mem[5530] <= 30'b000000010000000000101010000000
                ;mem[5531] <= 30'b000000010000000000101010010000
                ;mem[5532] <= 30'b000000010000000000101010100000
                ;mem[5533] <= 30'b000000010000000000101010110000
                ;mem[5534] <= 30'b000000010000000000101011000000
                ;mem[5535] <= 30'b000000010000000000110000100000
                ;mem[5536] <= 30'b000000010000000000110000110000
                ;mem[5537] <= 30'b000000010000000000110001110000
                ;mem[5538] <= 30'b000000010000000000110010000000
                ;mem[5539] <= 30'b000000010000000000110111010000
                ;mem[5540] <= 30'b000000010000000000110111100000
                ;mem[5541] <= 30'b000000010000000000111110010000
                ;mem[5542] <= 30'b000000010000000000111110100000
                ;mem[5543] <= 30'b000000000000000001000100100000
                ;mem[5544] <= 30'b000000000000000001000100110000
                ;mem[5545] <= 30'b000000000000000001000101110000
                ;mem[5546] <= 30'b000000000000000001000110000000
                ;mem[5547] <= 30'b000000000000000001001011010000
                ;mem[5548] <= 30'b000000000000000001001011100000
                ;mem[5549] <= 30'b000000000000000001010010010000
                ;mem[5550] <= 30'b000000000000000001010010100000
                ;mem[5551] <= 30'b000000000000000001011001000000
                ;mem[5552] <= 30'b000000000000000001011001010000
                ;mem[5553] <= 30'b000000000000000001100000000000
                ;mem[5554] <= 30'b000000000000000001100110110000
                ;mem[5555] <= 30'b000000000000000001100111000000
                ;mem[5556] <= 30'b000000000000000001101101110000
                ;mem[5557] <= 30'b000000000000000001110100110000
                ;mem[5558] <= 30'b000000000000000000101100010000
                ;mem[5559] <= 30'b000000000000000000101100100000
                ;mem[5560] <= 30'b000000000000000000101110100000
                ;mem[5561] <= 30'b000000000000000000101110110000
                ;mem[5562] <= 30'b000000000000000000110011000000
                ;mem[5563] <= 30'b000000000000000000110011010000
                ;mem[5564] <= 30'b000000000000000000110011100000
                ;mem[5565] <= 30'b000000000000000000110101100000
                ;mem[5566] <= 30'b000000000000000000110101110000
                ;mem[5567] <= 30'b000000000000000000111010000000
                ;mem[5568] <= 30'b000000000000000000111010010000
                ;mem[5569] <= 30'b000000000000000000111100010000
                ;mem[5570] <= 30'b000000000000000000111100100000
                ;mem[5571] <= 30'b000000000000000000111100110000
                ;mem[5572] <= 30'b000000001000000000000000010000
                ;mem[5573] <= 30'b000000001000000000000000100000
                ;mem[5574] <= 30'b000000001000000000000010100000
                ;mem[5575] <= 30'b000000001000000000000010110000
                ;mem[5576] <= 30'b000000001000000000000111000000
                ;mem[5577] <= 30'b000000001000000000000111010000
                ;mem[5578] <= 30'b000000001000000000000111100000
                ;mem[5579] <= 30'b000000001000000000001001100000
                ;mem[5580] <= 30'b000000001000000000001001110000
                ;mem[5581] <= 30'b000000001000000000001110000000
                ;mem[5582] <= 30'b000000001000000000001110010000
                ;mem[5583] <= 30'b000000001000000000010000010000
                ;mem[5584] <= 30'b000000001000000000010000100000
                ;mem[5585] <= 30'b000000001000000000010000110000
                ;mem[5586] <= 30'b000000001000000000010101000000
                ;mem[5587] <= 30'b000000001000000000010101010000
                ;mem[5588] <= 30'b000000001000000000010111010000
                ;mem[5589] <= 30'b000000001000000000010111100000
                ;mem[5590] <= 30'b000000001000000000010111110000
                ;mem[5591] <= 30'b000000001000000000011100000000
                ;mem[5592] <= 30'b000000001000000000011100010000
                ;mem[5593] <= 30'b000000001000000000011110000000
                ;mem[5594] <= 30'b000000001000000000011110010000
                ;mem[5595] <= 30'b000000001000000000011110100000
                ;mem[5596] <= 30'b000000001000000000011110110000
                ;mem[5597] <= 30'b000000001000000000100011000000
                ;mem[5598] <= 30'b000000001000000000100011010000
                ;mem[5599] <= 30'b000000001000000000100100110000
                ;mem[5600] <= 30'b000000001000000000100101000000
                ;mem[5601] <= 30'b000000001000000000100101010000
                ;mem[5602] <= 30'b000000001000000000100101100000
                ;mem[5603] <= 30'b000000001000000000101001110000
                ;mem[5604] <= 30'b000000001000000000101010000000
                ;mem[5605] <= 30'b000000001000000000101010010000
                ;mem[5606] <= 30'b000000001000000000101011110000
                ;mem[5607] <= 30'b000000001000000000101100000000
                ;mem[5608] <= 30'b000000001000000000101100010000
                ;mem[5609] <= 30'b000000001000000000101100100000
                ;mem[5610] <= 30'b000000001000000000110000110000
                ;mem[5611] <= 30'b000000001000000000110001000000
                ;mem[5612] <= 30'b000000001000000000110001010000
                ;mem[5613] <= 30'b000000001000000000110010100000
                ;mem[5614] <= 30'b000000001000000000110010110000
                ;mem[5615] <= 30'b000000001000000000110011000000
                ;mem[5616] <= 30'b000000001000000000110011010000
                ;mem[5617] <= 30'b000000001000000000110011100000
                ;mem[5618] <= 30'b000000001000000000111000000000
                ;mem[5619] <= 30'b000000001000000000111000010000
                ;mem[5620] <= 30'b000000001000000000111001010000
                ;mem[5621] <= 30'b000000001000000000111001100000
                ;mem[5622] <= 30'b000000001000000000111001110000
                ;mem[5623] <= 30'b000000001000000000111010000000
                ;mem[5624] <= 30'b000000001000000000111010010000
                ;mem[5625] <= 30'b000000001000000000111010100000
                ;mem[5626] <= 30'b000000001000000000111111000000
                ;mem[5627] <= 30'b000000001000000000111111010000
                ;mem[5628] <= 30'b000000001000000000111111100000
                ;mem[5629] <= 30'b000000010000000000000000000000
                ;mem[5630] <= 30'b000000010000000000000000010000
                ;mem[5631] <= 30'b000000010000000000000000100000
                ;mem[5632] <= 30'b000000010000000000000100110000
                ;mem[5633] <= 30'b000000010000000000000101000000
                ;mem[5634] <= 30'b000000010000000000000101010000
                ;mem[5635] <= 30'b000000010000000000000110100000
                ;mem[5636] <= 30'b000000010000000000000110110000
                ;mem[5637] <= 30'b000000010000000000000111000000
                ;mem[5638] <= 30'b000000010000000000000111010000
                ;mem[5639] <= 30'b000000010000000000000111100000
                ;mem[5640] <= 30'b000000010000000000001100000000
                ;mem[5641] <= 30'b000000010000000000001100010000
                ;mem[5642] <= 30'b000000010000000000001101010000
                ;mem[5643] <= 30'b000000010000000000001101100000
                ;mem[5644] <= 30'b000000010000000000001101110000
                ;mem[5645] <= 30'b000000010000000000001110000000
                ;mem[5646] <= 30'b000000010000000000001110010000
                ;mem[5647] <= 30'b000000010000000000001110100000
                ;mem[5648] <= 30'b000000010000000000010011000000
                ;mem[5649] <= 30'b000000010000000000010011010000
                ;mem[5650] <= 30'b000000010000000000010011100000
                ;mem[5651] <= 30'b000000010000000000010100000000
                ;mem[5652] <= 30'b000000010000000000010100010000
                ;mem[5653] <= 30'b000000010000000000010100100000
                ;mem[5654] <= 30'b000000010000000000010100110000
                ;mem[5655] <= 30'b000000010000000000010101000000
                ;mem[5656] <= 30'b000000010000000000010101010000
                ;mem[5657] <= 30'b000000010000000000011010010000
                ;mem[5658] <= 30'b000000010000000000011010100000
                ;mem[5659] <= 30'b000000010000000000011010110000
                ;mem[5660] <= 30'b000000010000000000011011000000
                ;mem[5661] <= 30'b000000010000000000011011010000
                ;mem[5662] <= 30'b000000010000000000011011100000
                ;mem[5663] <= 30'b000000010000000000011011110000
                ;mem[5664] <= 30'b000000010000000000011100000000
                ;mem[5665] <= 30'b000000010000000000011100010000
                ;mem[5666] <= 30'b000000010000000000100001110000
                ;mem[5667] <= 30'b000000010000000000100010000000
                ;mem[5668] <= 30'b000000010000000000100010110000
                ;mem[5669] <= 30'b000000010000000000100011000000
                ;mem[5670] <= 30'b000000010000000000100011010000
                ;mem[5671] <= 30'b000000010000000000101001100000
                ;mem[5672] <= 30'b000000010000000000101001110000
                ;mem[5673] <= 30'b000000010000000000101010000000
                ;mem[5674] <= 30'b000000010000000000101010010000
                ;mem[5675] <= 30'b000000010000000000110000100000
                ;mem[5676] <= 30'b000000010000000000110000110000
                ;mem[5677] <= 30'b000000010000000000110001000000
                ;mem[5678] <= 30'b000000010000000000110111100000
                ;mem[5679] <= 30'b000000010000000000110111110000
                ;mem[5680] <= 30'b000000010000000000111000000000
                ;mem[5681] <= 30'b000000010000000000111110100000
                ;mem[5682] <= 30'b000000010000000000111110110000
                ;mem[5683] <= 30'b000000000000000001000100100000
                ;mem[5684] <= 30'b000000000000000001000100110000
                ;mem[5685] <= 30'b000000000000000001000101000000
                ;mem[5686] <= 30'b000000000000000001001011100000
                ;mem[5687] <= 30'b000000000000000001001011110000
                ;mem[5688] <= 30'b000000000000000001001100000000
                ;mem[5689] <= 30'b000000000000000001010010100000
                ;mem[5690] <= 30'b000000000000000001010010110000
                ;mem[5691] <= 30'b000000000000000001011001100000
                ;mem[5692] <= 30'b000000000000000001011001110000
                ;mem[5693] <= 30'b000000000000000001100000100000
                ;mem[5694] <= 30'b000000000000000001100000110000
                ;mem[5695] <= 30'b000000000000000001100111100000
                ;mem[5696] <= 30'b000000000000000001100111110000
                ;mem[5697] <= 30'b000000000000000001101110110000
                ;mem[5698] <= 30'b000000000000000000100110110000
                ;mem[5699] <= 30'b000000000000000000100111000000
                ;mem[5700] <= 30'b000000000000000000100111010000
                ;mem[5701] <= 30'b000000000000000000101110000000
                ;mem[5702] <= 30'b000000000000000000101110010000
                ;mem[5703] <= 30'b000000000000000000110101000000
                ;mem[5704] <= 30'b000000000000000000110101010000
                ;mem[5705] <= 30'b000000000000000000111100000000
                ;mem[5706] <= 30'b000000000000000000111100010000
                ;mem[5707] <= 30'b000000001000000000000010000000
                ;mem[5708] <= 30'b000000001000000000000010010000
                ;mem[5709] <= 30'b000000001000000000001001000000
                ;mem[5710] <= 30'b000000001000000000001001010000
                ;mem[5711] <= 30'b000000001000000000010000000000
                ;mem[5712] <= 30'b000000001000000000010000010000
                ;mem[5713] <= 30'b000000001000000000010111000000
                ;mem[5714] <= 30'b000000001000000000011101110000
                ;mem[5715] <= 30'b000000001000000000011110000000
                ;mem[5716] <= 30'b000000001000000000100100100000
                ;mem[5717] <= 30'b000000001000000000100100110000
                ;mem[5718] <= 30'b000000001000000000101011010000
                ;mem[5719] <= 30'b000000001000000000101011100000
                ;mem[5720] <= 30'b000000001000000000101011110000
                ;mem[5721] <= 30'b000000001000000000110010010000
                ;mem[5722] <= 30'b000000001000000000110010100000
                ;mem[5723] <= 30'b000000001000000000111001000000
                ;mem[5724] <= 30'b000000001000000000111001010000
                ;mem[5725] <= 30'b000000001000000000111111110000
                ;mem[5726] <= 30'b000000010000000000000110010000
                ;mem[5727] <= 30'b000000010000000000000110100000
                ;mem[5728] <= 30'b000000010000000000001101000000
                ;mem[5729] <= 30'b000000010000000000001101010000
                ;mem[5730] <= 30'b000000010000000000010011110000
                ;mem[5731] <= 30'b000000010000000000010100000000
                ;mem[5732] <= 30'b000000010000000000010110100000
                ;mem[5733] <= 30'b000000010000000000010110110000
                ;mem[5734] <= 30'b000000010000000000011010110000
                ;mem[5735] <= 30'b000000010000000000011011000000
                ;mem[5736] <= 30'b000000010000000000011011010000
                ;mem[5737] <= 30'b000000010000000000011011100000
                ;mem[5738] <= 30'b000000010000000000011011110000
                ;mem[5739] <= 30'b000000010000000000011100000000
                ;mem[5740] <= 30'b000000010000000000011100010000
                ;mem[5741] <= 30'b000000010000000000011100100000
                ;mem[5742] <= 30'b000000010000000000011100110000
                ;mem[5743] <= 30'b000000010000000000011101000000
                ;mem[5744] <= 30'b000000010000000000011101010000
                ;mem[5745] <= 30'b000000010000000000011101100000
                ;mem[5746] <= 30'b000000010000000000011101110000
                ;mem[5747] <= 30'b000000010000000000100001010000
                ;mem[5748] <= 30'b000000010000000000100001100000
                ;mem[5749] <= 30'b000000010000000000100001110000
                ;mem[5750] <= 30'b000000010000000000100010000000
                ;mem[5751] <= 30'b000000010000000000100010010000
                ;mem[5752] <= 30'b000000010000000000100010100000
                ;mem[5753] <= 30'b000000010000000000100100110000
                ;mem[5754] <= 30'b000000010000000000100101000000
                ;mem[5755] <= 30'b000000010000000000100111110000
                ;mem[5756] <= 30'b000000010000000000101000000000
                ;mem[5757] <= 30'b000000010000000000101000010000
                ;mem[5758] <= 30'b000000010000000000101000100000
                ;mem[5759] <= 30'b000000010000000000101000110000
                ;mem[5760] <= 30'b000000010000000000101110010000
                ;mem[5761] <= 30'b000000010000000000101110100000
                ;mem[5762] <= 30'b000000010000000000101110110000
                ;mem[5763] <= 30'b000000010000000000101111000000
                ;mem[5764] <= 30'b000000010000000000101111010000
                ;mem[5765] <= 30'b000000010000000000110101010000
                ;mem[5766] <= 30'b000000010000000000110101100000
                ;mem[5767] <= 30'b000000010000000000110101110000
                ;mem[5768] <= 30'b000000010000000000110110000000
                ;mem[5769] <= 30'b000000000000000001000010010000
                ;mem[5770] <= 30'b000000000000000001000010100000
                ;mem[5771] <= 30'b000000000000000001000010110000
                ;mem[5772] <= 30'b000000000000000001000011000000
                ;mem[5773] <= 30'b000000000000000001000011010000
                ;mem[5774] <= 30'b000000000000000001001001010000
                ;mem[5775] <= 30'b000000000000000001001001100000
                ;mem[5776] <= 30'b000000000000000001001001110000
                ;mem[5777] <= 30'b000000000000000001001010000000
                ;mem[5778] <= 30'b000000000000000000011110100000
                ;mem[5779] <= 30'b000000000000000000011110110000
                ;mem[5780] <= 30'b000000000000000000011111000000
                ;mem[5781] <= 30'b000000000000000000011111010000
                ;mem[5782] <= 30'b000000000000000000100101010000
                ;mem[5783] <= 30'b000000000000000000100101100000
                ;mem[5784] <= 30'b000000000000000000100101110000
                ;mem[5785] <= 30'b000000000000000000100110000000
                ;mem[5786] <= 30'b000000000000000000100110010000
                ;mem[5787] <= 30'b000000000000000000101100000000
                ;mem[5788] <= 30'b000000000000000000101100010000
                ;mem[5789] <= 30'b000000000000000000101100100000
                ;mem[5790] <= 30'b000000000000000000101100110000
                ;mem[5791] <= 30'b000000000000000000101101000000
                ;mem[5792] <= 30'b000000000000000000101101010000
                ;mem[5793] <= 30'b000000000000000000101101100000
                ;mem[5794] <= 30'b000000000000000000110011000000
                ;mem[5795] <= 30'b000000000000000000110100000000
                ;mem[5796] <= 30'b000000000000000000110100010000
                ;mem[5797] <= 30'b000000000000000000110100100000
                ;mem[5798] <= 30'b000000000000000000111011010000
                ;mem[5799] <= 30'b000000000000000000111011100000
                ;mem[5800] <= 30'b000000001000000000000000000000
                ;mem[5801] <= 30'b000000001000000000000000010000
                ;mem[5802] <= 30'b000000001000000000000000100000
                ;mem[5803] <= 30'b000000001000000000000000110000
                ;mem[5804] <= 30'b000000001000000000000001000000
                ;mem[5805] <= 30'b000000001000000000000001010000
                ;mem[5806] <= 30'b000000001000000000000001100000
                ;mem[5807] <= 30'b000000001000000000000111000000
                ;mem[5808] <= 30'b000000001000000000001000000000
                ;mem[5809] <= 30'b000000001000000000001000010000
                ;mem[5810] <= 30'b000000001000000000001000100000
                ;mem[5811] <= 30'b000000001000000000001111010000
                ;mem[5812] <= 30'b000000001000000000001111100000
                ;mem[5813] <= 30'b000000001000000000010110010000
                ;mem[5814] <= 30'b000000001000000000010110100000
                ;mem[5815] <= 30'b000000001000000000011101010000
                ;mem[5816] <= 30'b000000001000000000011101100000
                ;mem[5817] <= 30'b000000001000000000100100000000
                ;mem[5818] <= 30'b000000001000000000100100010000
                ;mem[5819] <= 30'b000000001000000000100100100000
                ;mem[5820] <= 30'b000000001000000000101011000000
                ;mem[5821] <= 30'b000000001000000000101011010000
                ;mem[5822] <= 30'b000000001000000000101011100000
                ;mem[5823] <= 30'b000000001000000000110010000000
                ;mem[5824] <= 30'b000000001000000000110010010000
                ;mem[5825] <= 30'b000000001000000000110010100000
                ;mem[5826] <= 30'b000000001000000000110010110000
                ;mem[5827] <= 30'b000000001000000000110011000000
                ;mem[5828] <= 30'b000000001000000000111001000000
                ;mem[5829] <= 30'b000000001000000000111001010000
                ;mem[5830] <= 30'b000000001000000000111001100000
                ;mem[5831] <= 30'b000000001000000000111001110000
                ;mem[5832] <= 30'b000000001000000000111010000000
                ;mem[5833] <= 30'b000000001000000000111010010000
                ;mem[5834] <= 30'b000000010000000000000110000000
                ;mem[5835] <= 30'b000000010000000000000110010000
                ;mem[5836] <= 30'b000000010000000000000110100000
                ;mem[5837] <= 30'b000000010000000000000110110000
                ;mem[5838] <= 30'b000000010000000000000111000000
                ;mem[5839] <= 30'b000000010000000000001101000000
                ;mem[5840] <= 30'b000000010000000000001101010000
                ;mem[5841] <= 30'b000000010000000000001101100000
                ;mem[5842] <= 30'b000000010000000000001101110000
                ;mem[5843] <= 30'b000000010000000000001110000000
                ;mem[5844] <= 30'b000000010000000000001110010000
                ;mem[5845] <= 30'b000000010000000000010100110000
                ;mem[5846] <= 30'b000000010000000000010101000000
                ;mem[5847] <= 30'b000000010000000000010101010000
                ;mem[5848] <= 30'b000000010000000000010101100000
                ;mem[5849] <= 30'b000000010000000000011100000000
                ;mem[5850] <= 30'b000000010000000000011100010000
                ;mem[5851] <= 30'b000000010000000000011100100000
                ;mem[5852] <= 30'b000000010000000000100011000000
                ;mem[5853] <= 30'b000000010000000000100011010000
                ;mem[5854] <= 30'b000000010000000000100011100000
                ;mem[5855] <= 30'b000000010000000000101001110000
                ;mem[5856] <= 30'b000000010000000000101010000000
                ;mem[5857] <= 30'b000000010000000000101010010000
                ;mem[5858] <= 30'b000000010000000000101010100000
                ;mem[5859] <= 30'b000000010000000000110000100000
                ;mem[5860] <= 30'b000000010000000000110000110000
                ;mem[5861] <= 30'b000000010000000000110001000000
                ;mem[5862] <= 30'b000000010000000000110001010000
                ;mem[5863] <= 30'b000000010000000000110111000000
                ;mem[5864] <= 30'b000000010000000000110111010000
                ;mem[5865] <= 30'b000000010000000000110111100000
                ;mem[5866] <= 30'b000000010000000000110111110000
                ;mem[5867] <= 30'b000000010000000000111000000000
                ;mem[5868] <= 30'b000000010000000000111101110000
                ;mem[5869] <= 30'b000000010000000000111110000000
                ;mem[5870] <= 30'b000000010000000000111110010000
                ;mem[5871] <= 30'b000000010000000000111110100000
                ;mem[5872] <= 30'b000000010000000000111110110000
                ;mem[5873] <= 30'b000000000000000001000100100000
                ;mem[5874] <= 30'b000000000000000001000100110000
                ;mem[5875] <= 30'b000000000000000001000101000000
                ;mem[5876] <= 30'b000000000000000001000101010000
                ;mem[5877] <= 30'b000000000000000001001011000000
                ;mem[5878] <= 30'b000000000000000001001011010000
                ;mem[5879] <= 30'b000000000000000001001011100000
                ;mem[5880] <= 30'b000000000000000001001011110000
                ;mem[5881] <= 30'b000000000000000001001100000000
                ;mem[5882] <= 30'b000000000000000001010001110000
                ;mem[5883] <= 30'b000000000000000001010010000000
                ;mem[5884] <= 30'b000000000000000001010010010000
                ;mem[5885] <= 30'b000000000000000001010010100000
                ;mem[5886] <= 30'b000000000000000001010010110000
                ;mem[5887] <= 30'b000000000000000001011000100000
                ;mem[5888] <= 30'b000000000000000001011000110000
                ;mem[5889] <= 30'b000000000000000001011001000000
                ;mem[5890] <= 30'b000000000000000001011001010000
                ;mem[5891] <= 30'b000000000000000001011001100000
                ;mem[5892] <= 30'b000000000000000001011111110000
                ;mem[5893] <= 30'b000000000000000001100000000000
                ;mem[5894] <= 30'b000000000000000000100110000000
                ;mem[5895] <= 30'b000000000000000000100110010000
                ;mem[5896] <= 30'b000000000000000000100110100000
                ;mem[5897] <= 30'b000000000000000000101101000000
                ;mem[5898] <= 30'b000000000000000000101101010000
                ;mem[5899] <= 30'b000000000000000000101101100000
                ;mem[5900] <= 30'b000000000000000000101101110000
                ;mem[5901] <= 30'b000000000000000000101110000000
                ;mem[5902] <= 30'b000000000000000000101110010000
                ;mem[5903] <= 30'b000000000000000000101110100000
                ;mem[5904] <= 30'b000000000000000000101110110000
                ;mem[5905] <= 30'b000000000000000000101111000000
                ;mem[5906] <= 30'b000000000000000000110100000000
                ;mem[5907] <= 30'b000000000000000000110110010000
                ;mem[5908] <= 30'b000000000000000000111011000000
                ;mem[5909] <= 30'b000000001000000000000001000000
                ;mem[5910] <= 30'b000000001000000000000001010000
                ;mem[5911] <= 30'b000000001000000000000001100000
                ;mem[5912] <= 30'b000000001000000000000001110000
                ;mem[5913] <= 30'b000000001000000000000010000000
                ;mem[5914] <= 30'b000000001000000000000010010000
                ;mem[5915] <= 30'b000000001000000000000010100000
                ;mem[5916] <= 30'b000000001000000000000010110000
                ;mem[5917] <= 30'b000000001000000000000011000000
                ;mem[5918] <= 30'b000000001000000000001000000000
                ;mem[5919] <= 30'b000000001000000000001010010000
                ;mem[5920] <= 30'b000000001000000000001111000000
                ;mem[5921] <= 30'b000000001000000000010110000000
                ;mem[5922] <= 30'b000000001000000000011101000000
                ;mem[5923] <= 30'b000000001000000000100011110000
                ;mem[5924] <= 30'b000000001000000000100100000000
                ;mem[5925] <= 30'b000000001000000000101010110000
                ;mem[5926] <= 30'b000000001000000000101011000000
                ;mem[5927] <= 30'b000000001000000000101011010000
                ;mem[5928] <= 30'b000000001000000000101011100000
                ;mem[5929] <= 30'b000000001000000000101011110000
                ;mem[5930] <= 30'b000000001000000000101100000000
                ;mem[5931] <= 30'b000000001000000000110001110000
                ;mem[5932] <= 30'b000000001000000000110010000000
                ;mem[5933] <= 30'b000000001000000000110010010000
                ;mem[5934] <= 30'b000000001000000000110010100000
                ;mem[5935] <= 30'b000000001000000000110010110000
                ;mem[5936] <= 30'b000000001000000000110011000000
                ;mem[5937] <= 30'b000000001000000000110011010000
                ;mem[5938] <= 30'b000000001000000000111000100000
                ;mem[5939] <= 30'b000000001000000000111000110000
                ;mem[5940] <= 30'b000000001000000000111001000000
                ;mem[5941] <= 30'b000000001000000000111010010000
                ;mem[5942] <= 30'b000000001000000000111010100000
                ;mem[5943] <= 30'b000000001000000000111111010000
                ;mem[5944] <= 30'b000000001000000000111111100000
                ;mem[5945] <= 30'b000000001000000000111111110000
                ;mem[5946] <= 30'b000000010000000000000000000000
                ;mem[5947] <= 30'b000000010000000000000101110000
                ;mem[5948] <= 30'b000000010000000000000110000000
                ;mem[5949] <= 30'b000000010000000000000110010000
                ;mem[5950] <= 30'b000000010000000000000110100000
                ;mem[5951] <= 30'b000000010000000000000110110000
                ;mem[5952] <= 30'b000000010000000000000111000000
                ;mem[5953] <= 30'b000000010000000000000111010000
                ;mem[5954] <= 30'b000000010000000000001100100000
                ;mem[5955] <= 30'b000000010000000000001100110000
                ;mem[5956] <= 30'b000000010000000000001101000000
                ;mem[5957] <= 30'b000000010000000000001110010000
                ;mem[5958] <= 30'b000000010000000000001110100000
                ;mem[5959] <= 30'b000000010000000000010011010000
                ;mem[5960] <= 30'b000000010000000000010011100000
                ;mem[5961] <= 30'b000000010000000000010011110000
                ;mem[5962] <= 30'b000000010000000000010101010000
                ;mem[5963] <= 30'b000000010000000000010101100000
                ;mem[5964] <= 30'b000000010000000000011010100000
                ;mem[5965] <= 30'b000000010000000000011100100000
                ;mem[5966] <= 30'b000000010000000000100011100000
                ;mem[5967] <= 30'b000000010000000000101000010000
                ;mem[5968] <= 30'b000000010000000000101010010000
                ;mem[5969] <= 30'b000000010000000000101010100000
                ;mem[5970] <= 30'b000000010000000000101111000000
                ;mem[5971] <= 30'b000000010000000000101111010000
                ;mem[5972] <= 30'b000000010000000000110001010000
                ;mem[5973] <= 30'b000000010000000000110001100000
                ;mem[5974] <= 30'b000000010000000000110110000000
                ;mem[5975] <= 30'b000000010000000000111000000000
                ;mem[5976] <= 30'b000000010000000000111000010000
                ;mem[5977] <= 30'b000000010000000000111000100000
                ;mem[5978] <= 30'b000000010000000000111101000000
                ;mem[5979] <= 30'b000000010000000000111110110000
                ;mem[5980] <= 30'b000000010000000000111111000000
                ;mem[5981] <= 30'b000000010000000000111111010000
                ;mem[5982] <= 30'b000000000000000001000011000000
                ;mem[5983] <= 30'b000000000000000001000011010000
                ;mem[5984] <= 30'b000000000000000001000101010000
                ;mem[5985] <= 30'b000000000000000001000101100000
                ;mem[5986] <= 30'b000000000000000001001010000000
                ;mem[5987] <= 30'b000000000000000001001100000000
                ;mem[5988] <= 30'b000000000000000001001100010000
                ;mem[5989] <= 30'b000000000000000001001100100000
                ;mem[5990] <= 30'b000000000000000001010001000000
                ;mem[5991] <= 30'b000000000000000001010010110000
                ;mem[5992] <= 30'b000000000000000001010011000000
                ;mem[5993] <= 30'b000000000000000001010011010000
                ;mem[5994] <= 30'b000000000000000001011000000000
                ;mem[5995] <= 30'b000000000000000001011000010000
                ;mem[5996] <= 30'b000000000000000001011001010000
                ;mem[5997] <= 30'b000000000000000001011001100000
                ;mem[5998] <= 30'b000000000000000001011001110000
                ;mem[5999] <= 30'b000000000000000001011010000000
                ;mem[6000] <= 30'b000000000000000001011111010000
                ;mem[6001] <= 30'b000000000000000001011111100000
                ;mem[6002] <= 30'b000000000000000001011111110000
                ;mem[6003] <= 30'b000000000000000001100000000000
                ;mem[6004] <= 30'b000000000000000001100000010000
                ;mem[6005] <= 30'b000000000000000001100000100000
                ;mem[6006] <= 30'b000000000000000001100110100000
                ;mem[6007] <= 30'b000000000000000001100110110000
                ;mem[6008] <= 30'b000000000000000000011110100000
                ;mem[6009] <= 30'b000000000000000000011110110000
                ;mem[6010] <= 30'b000000000000000000011111000000
                ;mem[6011] <= 30'b000000000000000000100101100000
                ;mem[6012] <= 30'b000000000000000000100101110000
                ;mem[6013] <= 30'b000000000000000000100110000000
                ;mem[6014] <= 30'b000000000000000000101100100000
                ;mem[6015] <= 30'b000000000000000000101100110000
                ;mem[6016] <= 30'b000000000000000000101101000000
                ;mem[6017] <= 30'b000000000000000000101101010000
                ;mem[6018] <= 30'b000000000000000000110011100000
                ;mem[6019] <= 30'b000000000000000000110011110000
                ;mem[6020] <= 30'b000000000000000000110100000000
                ;mem[6021] <= 30'b000000000000000000110100010000
                ;mem[6022] <= 30'b000000000000000000111010110000
                ;mem[6023] <= 30'b000000000000000000111011000000
                ;mem[6024] <= 30'b000000000000000000111011010000
                ;mem[6025] <= 30'b000000000000000000111011100000
                ;mem[6026] <= 30'b000000001000000000000000100000
                ;mem[6027] <= 30'b000000001000000000000000110000
                ;mem[6028] <= 30'b000000001000000000000001000000
                ;mem[6029] <= 30'b000000001000000000000001010000
                ;mem[6030] <= 30'b000000001000000000000111100000
                ;mem[6031] <= 30'b000000001000000000000111110000
                ;mem[6032] <= 30'b000000001000000000001000000000
                ;mem[6033] <= 30'b000000001000000000001000010000
                ;mem[6034] <= 30'b000000001000000000001110110000
                ;mem[6035] <= 30'b000000001000000000001111000000
                ;mem[6036] <= 30'b000000001000000000001111010000
                ;mem[6037] <= 30'b000000001000000000001111100000
                ;mem[6038] <= 30'b000000001000000000010101110000
                ;mem[6039] <= 30'b000000001000000000010110000000
                ;mem[6040] <= 30'b000000001000000000010110010000
                ;mem[6041] <= 30'b000000001000000000010110100000
                ;mem[6042] <= 30'b000000001000000000011101000000
                ;mem[6043] <= 30'b000000001000000000011101010000
                ;mem[6044] <= 30'b000000001000000000011101100000
                ;mem[6045] <= 30'b000000001000000000011101110000
                ;mem[6046] <= 30'b000000001000000000100100000000
                ;mem[6047] <= 30'b000000001000000000100100010000
                ;mem[6048] <= 30'b000000001000000000100100100000
                ;mem[6049] <= 30'b000000001000000000100100110000
                ;mem[6050] <= 30'b000000001000000000101011010000
                ;mem[6051] <= 30'b000000001000000000101011100000
                ;mem[6052] <= 30'b000000001000000000101011110000
                ;mem[6053] <= 30'b000000001000000000110010010000
                ;mem[6054] <= 30'b000000001000000000110010100000
                ;mem[6055] <= 30'b000000001000000000110010110000
                ;mem[6056] <= 30'b000000001000000000110011000000
                ;mem[6057] <= 30'b000000001000000000111001010000
                ;mem[6058] <= 30'b000000001000000000111001100000
                ;mem[6059] <= 30'b000000001000000000111001110000
                ;mem[6060] <= 30'b000000001000000000111010000000
                ;mem[6061] <= 30'b000000010000000000000110010000
                ;mem[6062] <= 30'b000000010000000000000110100000
                ;mem[6063] <= 30'b000000010000000000000110110000
                ;mem[6064] <= 30'b000000010000000000000111000000
                ;mem[6065] <= 30'b000000010000000000001101010000
                ;mem[6066] <= 30'b000000010000000000001101100000
                ;mem[6067] <= 30'b000000010000000000001101110000
                ;mem[6068] <= 30'b000000010000000000001110000000
                ;mem[6069] <= 30'b000000010000000000010100010000
                ;mem[6070] <= 30'b000000010000000000010100100000
                ;mem[6071] <= 30'b000000010000000000010100110000
                ;mem[6072] <= 30'b000000010000000000010101000000
                ;mem[6073] <= 30'b000000010000000000011011100000
                ;mem[6074] <= 30'b000000010000000000011011110000
                ;mem[6075] <= 30'b000000010000000000011100000000
                ;mem[6076] <= 30'b000000010000000000011100010000
                ;mem[6077] <= 30'b000000010000000000100010100000
                ;mem[6078] <= 30'b000000010000000000100010110000
                ;mem[6079] <= 30'b000000010000000000100011000000
                ;mem[6080] <= 30'b000000010000000000100011010000
                ;mem[6081] <= 30'b000000010000000000101001110000
                ;mem[6082] <= 30'b000000010000000000101010000000
                ;mem[6083] <= 30'b000000010000000000101010010000
                ;mem[6084] <= 30'b000000010000000000101010100000
                ;mem[6085] <= 30'b000000010000000000110000110000
                ;mem[6086] <= 30'b000000010000000000110001000000
                ;mem[6087] <= 30'b000000010000000000110001010000
                ;mem[6088] <= 30'b000000010000000000110001100000
                ;mem[6089] <= 30'b000000010000000000110111110000
                ;mem[6090] <= 30'b000000010000000000111000000000
                ;mem[6091] <= 30'b000000010000000000111000010000
                ;mem[6092] <= 30'b000000010000000000111000100000
                ;mem[6093] <= 30'b000000010000000000111000110000
                ;mem[6094] <= 30'b000000010000000000111111000000
                ;mem[6095] <= 30'b000000010000000000111111010000
                ;mem[6096] <= 30'b000000010000000000111111100000
                ;mem[6097] <= 30'b000000010000000000111111110000
                ;mem[6098] <= 30'b000000000000000001000100110000
                ;mem[6099] <= 30'b000000000000000001000101000000
                ;mem[6100] <= 30'b000000000000000001000101010000
                ;mem[6101] <= 30'b000000000000000001000101100000
                ;mem[6102] <= 30'b000000000000000001001011110000
                ;mem[6103] <= 30'b000000000000000001001100000000
                ;mem[6104] <= 30'b000000000000000001001100010000
                ;mem[6105] <= 30'b000000000000000001001100100000
                ;mem[6106] <= 30'b000000000000000001001100110000
                ;mem[6107] <= 30'b000000000000000001010011000000
                ;mem[6108] <= 30'b000000000000000001010011010000
                ;mem[6109] <= 30'b000000000000000001010011100000
                ;mem[6110] <= 30'b000000000000000001010011110000
                ;mem[6111] <= 30'b000000000000000001011010000000
                ;mem[6112] <= 30'b000000000000000001011010010000
                ;mem[6113] <= 30'b000000000000000001011010100000
                ;mem[6114] <= 30'b000000000000000001100001010000
                ;mem[6115] <= 30'b000000000000000001100001100000
                ;mem[6116] <= 30'b000000000000000000010000100000
                ;mem[6117] <= 30'b000000000000000000010000110000
                ;mem[6118] <= 30'b000000000000000000010001000000
                ;mem[6119] <= 30'b000000000000000000010001010000
                ;mem[6120] <= 30'b000000000000000000010111010000
                ;mem[6121] <= 30'b000000000000000000011000010000
                ;mem[6122] <= 30'b000000000000000000011000100000
                ;mem[6123] <= 30'b000000000000000000011111110000
                ;mem[6124] <= 30'b000000000000000000100111000000
                ;mem[6125] <= 30'b000000000000000000101110000000
                ;mem[6126] <= 30'b000000000000000000101110010000
                ;mem[6127] <= 30'b000000000000000000110101010000
                ;mem[6128] <= 30'b000000000000000000111100010000
                ;mem[6129] <= 30'b000000001000000000000010000000
                ;mem[6130] <= 30'b000000001000000000000010010000
                ;mem[6131] <= 30'b000000001000000000001001010000
                ;mem[6132] <= 30'b000000001000000000010000010000
                ;mem[6133] <= 30'b000000001000000000010111010000
                ;mem[6134] <= 30'b000000001000000000010111100000
                ;mem[6135] <= 30'b000000001000000000011110010000
                ;mem[6136] <= 30'b000000001000000000011110100000
                ;mem[6137] <= 30'b000000001000000000100101010000
                ;mem[6138] <= 30'b000000001000000000100101100000
                ;mem[6139] <= 30'b000000001000000000101100010000
                ;mem[6140] <= 30'b000000001000000000110011010000
                ;mem[6141] <= 30'b000000001000000000111010000000
                ;mem[6142] <= 30'b000000001000000000111010010000
                ;mem[6143] <= 30'b000000001000000000111111010000
                ;mem[6144] <= 30'b000000001000000000111111100000
                ;mem[6145] <= 30'b000000001000000000111111110000
                ;mem[6146] <= 30'b000000010000000000000000010000
                ;mem[6147] <= 30'b000000010000000000000111010000
                ;mem[6148] <= 30'b000000010000000000001110000000
                ;mem[6149] <= 30'b000000010000000000001110010000
                ;mem[6150] <= 30'b000000010000000000010011010000
                ;mem[6151] <= 30'b000000010000000000010011100000
                ;mem[6152] <= 30'b000000010000000000010011110000
                ;mem[6153] <= 30'b000000010000000000010100000000
                ;mem[6154] <= 30'b000000010000000000010100010000
                ;mem[6155] <= 30'b000000010000000000010101000000
                ;mem[6156] <= 30'b000000010000000000011010000000
                ;mem[6157] <= 30'b000000010000000000011010010000
                ;mem[6158] <= 30'b000000010000000000011011100000
                ;mem[6159] <= 30'b000000010000000000011011110000
                ;mem[6160] <= 30'b000000010000000000011100000000
                ;mem[6161] <= 30'b000000010000000000100001000000
                ;mem[6162] <= 30'b000000010000000000100010110000
                ;mem[6163] <= 30'b000000010000000000100011000000
                ;mem[6164] <= 30'b000000010000000000101000000000
                ;mem[6165] <= 30'b000000010000000000101001100000
                ;mem[6166] <= 30'b000000010000000000101001110000
                ;mem[6167] <= 30'b000000010000000000101010000000
                ;mem[6168] <= 30'b000000010000000000101010010000
                ;mem[6169] <= 30'b000000010000000000101111000000
                ;mem[6170] <= 30'b000000010000000000110000010000
                ;mem[6171] <= 30'b000000010000000000110000100000
                ;mem[6172] <= 30'b000000010000000000110001010000
                ;mem[6173] <= 30'b000000010000000000110001100000
                ;mem[6174] <= 30'b000000010000000000110110000000
                ;mem[6175] <= 30'b000000010000000000110110010000
                ;mem[6176] <= 30'b000000010000000000110110100000
                ;mem[6177] <= 30'b000000010000000000110110110000
                ;mem[6178] <= 30'b000000010000000000110111000000
                ;mem[6179] <= 30'b000000010000000000110111010000
                ;mem[6180] <= 30'b000000010000000000111000100000
                ;mem[6181] <= 30'b000000010000000000111000110000
                ;mem[6182] <= 30'b000000010000000000111001000000
                ;mem[6183] <= 30'b000000010000000000111101010000
                ;mem[6184] <= 30'b000000010000000000111101100000
                ;mem[6185] <= 30'b000000000000000001000011000000
                ;mem[6186] <= 30'b000000000000000001000100010000
                ;mem[6187] <= 30'b000000000000000001000100100000
                ;mem[6188] <= 30'b000000000000000001000101010000
                ;mem[6189] <= 30'b000000000000000001000101100000
                ;mem[6190] <= 30'b000000000000000001001010000000
                ;mem[6191] <= 30'b000000000000000001001010010000
                ;mem[6192] <= 30'b000000000000000001001010100000
                ;mem[6193] <= 30'b000000000000000001001010110000
                ;mem[6194] <= 30'b000000000000000001001011000000
                ;mem[6195] <= 30'b000000000000000001001011010000
                ;mem[6196] <= 30'b000000000000000001001100100000
                ;mem[6197] <= 30'b000000000000000001001100110000
                ;mem[6198] <= 30'b000000000000000001001101000000
                ;mem[6199] <= 30'b000000000000000001010001010000
                ;mem[6200] <= 30'b000000000000000001010001100000
                ;mem[6201] <= 30'b000000000000000001010100000000
                ;mem[6202] <= 30'b000000000000000001010100010000
                ;mem[6203] <= 30'b000000000000000000101100110000
                ;mem[6204] <= 30'b000000000000000000101110110000
                ;mem[6205] <= 30'b000000000000000000101111000000
                ;mem[6206] <= 30'b000000000000000000110011100000
                ;mem[6207] <= 30'b000000000000000000110011110000
                ;mem[6208] <= 30'b000000000000000000110100000000
                ;mem[6209] <= 30'b000000000000000000110101100000
                ;mem[6210] <= 30'b000000000000000000110101110000
                ;mem[6211] <= 30'b000000000000000000110110000000
                ;mem[6212] <= 30'b000000000000000000111010010000
                ;mem[6213] <= 30'b000000000000000000111010100000
                ;mem[6214] <= 30'b000000000000000000111010110000
                ;mem[6215] <= 30'b000000000000000000111011000000
                ;mem[6216] <= 30'b000000000000000000111100010000
                ;mem[6217] <= 30'b000000000000000000111100100000
                ;mem[6218] <= 30'b000000000000000000111100110000
                ;mem[6219] <= 30'b000000000000000000111101000000
                ;mem[6220] <= 30'b000000001000000000000000110000
                ;mem[6221] <= 30'b000000001000000000000010110000
                ;mem[6222] <= 30'b000000001000000000000011000000
                ;mem[6223] <= 30'b000000001000000000000111100000
                ;mem[6224] <= 30'b000000001000000000000111110000
                ;mem[6225] <= 30'b000000001000000000001000000000
                ;mem[6226] <= 30'b000000001000000000001001100000
                ;mem[6227] <= 30'b000000001000000000001001110000
                ;mem[6228] <= 30'b000000001000000000001010000000
                ;mem[6229] <= 30'b000000001000000000001110010000
                ;mem[6230] <= 30'b000000001000000000001110100000
                ;mem[6231] <= 30'b000000001000000000001110110000
                ;mem[6232] <= 30'b000000001000000000001111000000
                ;mem[6233] <= 30'b000000001000000000010000010000
                ;mem[6234] <= 30'b000000001000000000010000100000
                ;mem[6235] <= 30'b000000001000000000010000110000
                ;mem[6236] <= 30'b000000001000000000010001000000
                ;mem[6237] <= 30'b000000001000000000010101000000
                ;mem[6238] <= 30'b000000001000000000010101010000
                ;mem[6239] <= 30'b000000001000000000010101100000
                ;mem[6240] <= 30'b000000001000000000010101110000
                ;mem[6241] <= 30'b000000001000000000010110000000
                ;mem[6242] <= 30'b000000001000000000010111010000
                ;mem[6243] <= 30'b000000001000000000010111100000
                ;mem[6244] <= 30'b000000001000000000010111110000
                ;mem[6245] <= 30'b000000001000000000011000000000
                ;mem[6246] <= 30'b000000001000000000011000010000
                ;mem[6247] <= 30'b000000001000000000011100000000
                ;mem[6248] <= 30'b000000001000000000011100010000
                ;mem[6249] <= 30'b000000001000000000011100100000
                ;mem[6250] <= 30'b000000001000000000011100110000
                ;mem[6251] <= 30'b000000001000000000011110010000
                ;mem[6252] <= 30'b000000001000000000011110100000
                ;mem[6253] <= 30'b000000001000000000011110110000
                ;mem[6254] <= 30'b000000001000000000011111000000
                ;mem[6255] <= 30'b000000001000000000100010110000
                ;mem[6256] <= 30'b000000001000000000100011000000
                ;mem[6257] <= 30'b000000001000000000100011010000
                ;mem[6258] <= 30'b000000001000000000100011100000
                ;mem[6259] <= 30'b000000001000000000100011110000
                ;mem[6260] <= 30'b000000001000000000100101000000
                ;mem[6261] <= 30'b000000001000000000100101010000
                ;mem[6262] <= 30'b000000001000000000100101100000
                ;mem[6263] <= 30'b000000001000000000100101110000
                ;mem[6264] <= 30'b000000001000000000100110000000
                ;mem[6265] <= 30'b000000001000000000101001110000
                ;mem[6266] <= 30'b000000001000000000101010000000
                ;mem[6267] <= 30'b000000001000000000101010010000
                ;mem[6268] <= 30'b000000001000000000101010100000
                ;mem[6269] <= 30'b000000001000000000101010110000
                ;mem[6270] <= 30'b000000001000000000101011100000
                ;mem[6271] <= 30'b000000001000000000101011110000
                ;mem[6272] <= 30'b000000001000000000101100000000
                ;mem[6273] <= 30'b000000001000000000101100010000
                ;mem[6274] <= 30'b000000001000000000101100100000
                ;mem[6275] <= 30'b000000001000000000101100110000
                ;mem[6276] <= 30'b000000001000000000101101000000
                ;mem[6277] <= 30'b000000001000000000110000100000
                ;mem[6278] <= 30'b000000001000000000110000110000
                ;mem[6279] <= 30'b000000001000000000110001000000
                ;mem[6280] <= 30'b000000001000000000110001010000
                ;mem[6281] <= 30'b000000001000000000110001100000
                ;mem[6282] <= 30'b000000001000000000110001110000
                ;mem[6283] <= 30'b000000001000000000110010000000
                ;mem[6284] <= 30'b000000001000000000110010010000
                ;mem[6285] <= 30'b000000001000000000110010100000
                ;mem[6286] <= 30'b000000001000000000110010110000
                ;mem[6287] <= 30'b000000001000000000110011000000
                ;mem[6288] <= 30'b000000001000000000110011010000
                ;mem[6289] <= 30'b000000001000000000110011100000
                ;mem[6290] <= 30'b000000001000000000110011110000
                ;mem[6291] <= 30'b000000001000000000110111110000
                ;mem[6292] <= 30'b000000001000000000111000000000
                ;mem[6293] <= 30'b000000001000000000111000010000
                ;mem[6294] <= 30'b000000001000000000111000100000
                ;mem[6295] <= 30'b000000001000000000111000110000
                ;mem[6296] <= 30'b000000001000000000111001000000
                ;mem[6297] <= 30'b000000001000000000111001010000
                ;mem[6298] <= 30'b000000001000000000111001100000
                ;mem[6299] <= 30'b000000001000000000111001110000
                ;mem[6300] <= 30'b000000001000000000111010000000
                ;mem[6301] <= 30'b000000001000000000111010010000
                ;mem[6302] <= 30'b000000001000000000111010100000
                ;mem[6303] <= 30'b000000001000000000111010110000
                ;mem[6304] <= 30'b000000001000000000111110110000
                ;mem[6305] <= 30'b000000001000000000111111000000
                ;mem[6306] <= 30'b000000001000000000111111010000
                ;mem[6307] <= 30'b000000001000000000111111100000
                ;mem[6308] <= 30'b000000001000000000111111110000
                ;mem[6309] <= 30'b000000010000000000000000000000
                ;mem[6310] <= 30'b000000010000000000000000010000
                ;mem[6311] <= 30'b000000010000000000000000100000
                ;mem[6312] <= 30'b000000010000000000000000110000
                ;mem[6313] <= 30'b000000010000000000000001000000
                ;mem[6314] <= 30'b000000010000000000000100100000
                ;mem[6315] <= 30'b000000010000000000000100110000
                ;mem[6316] <= 30'b000000010000000000000101000000
                ;mem[6317] <= 30'b000000010000000000000101010000
                ;mem[6318] <= 30'b000000010000000000000101100000
                ;mem[6319] <= 30'b000000010000000000000101110000
                ;mem[6320] <= 30'b000000010000000000000110000000
                ;mem[6321] <= 30'b000000010000000000000110010000
                ;mem[6322] <= 30'b000000010000000000000110100000
                ;mem[6323] <= 30'b000000010000000000000110110000
                ;mem[6324] <= 30'b000000010000000000000111000000
                ;mem[6325] <= 30'b000000010000000000000111010000
                ;mem[6326] <= 30'b000000010000000000000111100000
                ;mem[6327] <= 30'b000000010000000000000111110000
                ;mem[6328] <= 30'b000000010000000000001011110000
                ;mem[6329] <= 30'b000000010000000000001100000000
                ;mem[6330] <= 30'b000000010000000000001100010000
                ;mem[6331] <= 30'b000000010000000000001100100000
                ;mem[6332] <= 30'b000000010000000000001100110000
                ;mem[6333] <= 30'b000000010000000000001101000000
                ;mem[6334] <= 30'b000000010000000000001101010000
                ;mem[6335] <= 30'b000000010000000000001101100000
                ;mem[6336] <= 30'b000000010000000000001101110000
                ;mem[6337] <= 30'b000000010000000000001110000000
                ;mem[6338] <= 30'b000000010000000000001110010000
                ;mem[6339] <= 30'b000000010000000000001110100000
                ;mem[6340] <= 30'b000000010000000000001110110000
                ;mem[6341] <= 30'b000000010000000000010010110000
                ;mem[6342] <= 30'b000000010000000000010011000000
                ;mem[6343] <= 30'b000000010000000000010011010000
                ;mem[6344] <= 30'b000000010000000000010011100000
                ;mem[6345] <= 30'b000000010000000000010011110000
                ;mem[6346] <= 30'b000000010000000000010100000000
                ;mem[6347] <= 30'b000000010000000000010100010000
                ;mem[6348] <= 30'b000000010000000000010100100000
                ;mem[6349] <= 30'b000000010000000000010100110000
                ;mem[6350] <= 30'b000000010000000000010101000000
                ;mem[6351] <= 30'b000000010000000000010101010000
                ;mem[6352] <= 30'b000000010000000000010101100000
                ;mem[6353] <= 30'b000000010000000000010101110000
                ;mem[6354] <= 30'b000000010000000000011001110000
                ;mem[6355] <= 30'b000000010000000000011010000000
                ;mem[6356] <= 30'b000000010000000000011010010000
                ;mem[6357] <= 30'b000000010000000000011010100000
                ;mem[6358] <= 30'b000000010000000000011010110000
                ;mem[6359] <= 30'b000000010000000000011011000000
                ;mem[6360] <= 30'b000000010000000000011011010000
                ;mem[6361] <= 30'b000000010000000000011011100000
                ;mem[6362] <= 30'b000000010000000000011011110000
                ;mem[6363] <= 30'b000000010000000000011100000000
                ;mem[6364] <= 30'b000000010000000000011100010000
                ;mem[6365] <= 30'b000000010000000000011100100000
                ;mem[6366] <= 30'b000000010000000000011100110000
                ;mem[6367] <= 30'b000000010000000000100010110000
                ;mem[6368] <= 30'b000000010000000000100011000000
                ;mem[6369] <= 30'b000000010000000000100011010000
                ;mem[6370] <= 30'b000000010000000000100011100000
                ;mem[6371] <= 30'b000000010000000000101001110000
                ;mem[6372] <= 30'b000000010000000000101010000000
                ;mem[6373] <= 30'b000000010000000000101010010000
                ;mem[6374] <= 30'b000000010000000000101010100000
                ;mem[6375] <= 30'b000000010000000000110000110000
                ;mem[6376] <= 30'b000000010000000000110001000000
                ;mem[6377] <= 30'b000000010000000000110001010000
                ;mem[6378] <= 30'b000000010000000000110001100000
                ;mem[6379] <= 30'b000000010000000000110001110000
                ;mem[6380] <= 30'b000000010000000000110111110000
                ;mem[6381] <= 30'b000000010000000000111000000000
                ;mem[6382] <= 30'b000000010000000000111000010000
                ;mem[6383] <= 30'b000000010000000000111000100000
                ;mem[6384] <= 30'b000000010000000000111000110000
                ;mem[6385] <= 30'b000000010000000000111110100000
                ;mem[6386] <= 30'b000000010000000000111110110000
                ;mem[6387] <= 30'b000000010000000000111111000000
                ;mem[6388] <= 30'b000000010000000000111111010000
                ;mem[6389] <= 30'b000000010000000000111111100000
                ;mem[6390] <= 30'b000000000000000001000100110000
                ;mem[6391] <= 30'b000000000000000001000101000000
                ;mem[6392] <= 30'b000000000000000001000101010000
                ;mem[6393] <= 30'b000000000000000001000101100000
                ;mem[6394] <= 30'b000000000000000001000101110000
                ;mem[6395] <= 30'b000000000000000001001011110000
                ;mem[6396] <= 30'b000000000000000001001100000000
                ;mem[6397] <= 30'b000000000000000001001100010000
                ;mem[6398] <= 30'b000000000000000001001100100000
                ;mem[6399] <= 30'b000000000000000001001100110000
                ;mem[6400] <= 30'b000000000000000001010010100000
                ;mem[6401] <= 30'b000000000000000001010010110000
                ;mem[6402] <= 30'b000000000000000001010011000000
                ;mem[6403] <= 30'b000000000000000001010011010000
                ;mem[6404] <= 30'b000000000000000001010011100000
                ;mem[6405] <= 30'b000000000000000001011001100000
                ;mem[6406] <= 30'b000000000000000001011001110000
                ;mem[6407] <= 30'b000000000000000001011010000000
                ;mem[6408] <= 30'b000000000000000001011010010000
                ;mem[6409] <= 30'b000000000000000001011010100000
                ;mem[6410] <= 30'b000000000000000001100000100000
                ;mem[6411] <= 30'b000000000000000001100000110000
                ;mem[6412] <= 30'b000000000000000001100001000000
                ;mem[6413] <= 30'b000000000000000001100001010000
                ;mem[6414] <= 30'b000000000000000001100001100000
                ;mem[6415] <= 30'b000000000000000001100111100000
                ;mem[6416] <= 30'b000000000000000001100111110000
                ;mem[6417] <= 30'b000000000000000001101000000000
                ;mem[6418] <= 30'b000000000000000001101000010000
                ;mem[6419] <= 30'b000000000000000001101110100000
                ;mem[6420] <= 30'b000000000000000001101110110000
                ;mem[6421] <= 30'b000000000000000001101111000000
                ;mem[6422] <= 30'b000000000000000000100101000000
                ;mem[6423] <= 30'b000000000000000000101011110000
                ;mem[6424] <= 30'b000000000000000000101100000000
                ;mem[6425] <= 30'b000000000000000000101110100000
                ;mem[6426] <= 30'b000000000000000000110010110000
                ;mem[6427] <= 30'b000000000000000000110011000000
                ;mem[6428] <= 30'b000000000000000000110101100000
                ;mem[6429] <= 30'b000000000000000000110101110000
                ;mem[6430] <= 30'b000000000000000000111001110000
                ;mem[6431] <= 30'b000000000000000000111010000000
                ;mem[6432] <= 30'b000000000000000000111100100000
                ;mem[6433] <= 30'b000000000000000000111100110000
                ;mem[6434] <= 30'b000000001000000000000000000000
                ;mem[6435] <= 30'b000000001000000000000010100000
                ;mem[6436] <= 30'b000000001000000000000110110000
                ;mem[6437] <= 30'b000000001000000000000111000000
                ;mem[6438] <= 30'b000000001000000000001001100000
                ;mem[6439] <= 30'b000000001000000000001001110000
                ;mem[6440] <= 30'b000000001000000000001101110000
                ;mem[6441] <= 30'b000000001000000000001110000000
                ;mem[6442] <= 30'b000000001000000000010000100000
                ;mem[6443] <= 30'b000000001000000000010000110000
                ;mem[6444] <= 30'b000000001000000000010100110000
                ;mem[6445] <= 30'b000000001000000000010101000000
                ;mem[6446] <= 30'b000000001000000000010111100000
                ;mem[6447] <= 30'b000000001000000000010111110000
                ;mem[6448] <= 30'b000000001000000000011011110000
                ;mem[6449] <= 30'b000000001000000000011100000000
                ;mem[6450] <= 30'b000000001000000000011110100000
                ;mem[6451] <= 30'b000000001000000000011110110000
                ;mem[6452] <= 30'b000000001000000000100010110000
                ;mem[6453] <= 30'b000000001000000000100011000000
                ;mem[6454] <= 30'b000000001000000000100101100000
                ;mem[6455] <= 30'b000000001000000000100101110000
                ;mem[6456] <= 30'b000000001000000000100110100000
                ;mem[6457] <= 30'b000000001000000000101001110000
                ;mem[6458] <= 30'b000000001000000000101010000000
                ;mem[6459] <= 30'b000000001000000000101100100000
                ;mem[6460] <= 30'b000000001000000000101100110000
                ;mem[6461] <= 30'b000000001000000000101101010000
                ;mem[6462] <= 30'b000000001000000000101101100000
                ;mem[6463] <= 30'b000000001000000000110000110000
                ;mem[6464] <= 30'b000000001000000000110001000000
                ;mem[6465] <= 30'b000000001000000000110011010000
                ;mem[6466] <= 30'b000000001000000000110011100000
                ;mem[6467] <= 30'b000000001000000000110011110000
                ;mem[6468] <= 30'b000000001000000000110100000000
                ;mem[6469] <= 30'b000000001000000000110100010000
                ;mem[6470] <= 30'b000000001000000000110111110000
                ;mem[6471] <= 30'b000000001000000000111000000000
                ;mem[6472] <= 30'b000000001000000000111010010000
                ;mem[6473] <= 30'b000000001000000000111010100000
                ;mem[6474] <= 30'b000000001000000000111010110000
                ;mem[6475] <= 30'b000000001000000000111011000000
                ;mem[6476] <= 30'b000000001000000000111110110000
                ;mem[6477] <= 30'b000000001000000000111111000000
                ;mem[6478] <= 30'b000000001000000000111111010000
                ;mem[6479] <= 30'b000000001000000000111111100000
                ;mem[6480] <= 30'b000000010000000000000000100000
                ;mem[6481] <= 30'b000000010000000000000000110000
                ;mem[6482] <= 30'b000000010000000000000001010000
                ;mem[6483] <= 30'b000000010000000000000001100000
                ;mem[6484] <= 30'b000000010000000000000100110000
                ;mem[6485] <= 30'b000000010000000000000101000000
                ;mem[6486] <= 30'b000000010000000000000111010000
                ;mem[6487] <= 30'b000000010000000000000111100000
                ;mem[6488] <= 30'b000000010000000000000111110000
                ;mem[6489] <= 30'b000000010000000000001000000000
                ;mem[6490] <= 30'b000000010000000000001000010000
                ;mem[6491] <= 30'b000000010000000000001011110000
                ;mem[6492] <= 30'b000000010000000000001100000000
                ;mem[6493] <= 30'b000000010000000000001110010000
                ;mem[6494] <= 30'b000000010000000000001110100000
                ;mem[6495] <= 30'b000000010000000000001110110000
                ;mem[6496] <= 30'b000000010000000000001111000000
                ;mem[6497] <= 30'b000000010000000000010010110000
                ;mem[6498] <= 30'b000000010000000000010011000000
                ;mem[6499] <= 30'b000000010000000000010011010000
                ;mem[6500] <= 30'b000000010000000000010011100000
                ;mem[6501] <= 30'b000000010000000000010100100000
                ;mem[6502] <= 30'b000000010000000000010100110000
                ;mem[6503] <= 30'b000000010000000000010101000000
                ;mem[6504] <= 30'b000000010000000000010101010000
                ;mem[6505] <= 30'b000000010000000000010101100000
                ;mem[6506] <= 30'b000000010000000000010101110000
                ;mem[6507] <= 30'b000000010000000000011010000000
                ;mem[6508] <= 30'b000000010000000000011010010000
                ;mem[6509] <= 30'b000000010000000000011010100000
                ;mem[6510] <= 30'b000000010000000000011010110000
                ;mem[6511] <= 30'b000000010000000000011011000000
                ;mem[6512] <= 30'b000000010000000000011011010000
                ;mem[6513] <= 30'b000000010000000000011011100000
                ;mem[6514] <= 30'b000000010000000000011011110000
                ;mem[6515] <= 30'b000000010000000000011100000000
                ;mem[6516] <= 30'b000000010000000000011100010000
                ;mem[6517] <= 30'b000000010000000000011100100000
                ;mem[6518] <= 30'b000000010000000000011100110000
                ;mem[6519] <= 30'b000000010000000000100001010000
                ;mem[6520] <= 30'b000000010000000000100001100000
                ;mem[6521] <= 30'b000000010000000000100001110000
                ;mem[6522] <= 30'b000000010000000000100010000000
                ;mem[6523] <= 30'b000000010000000000100010010000
                ;mem[6524] <= 30'b000000010000000000100010100000
                ;mem[6525] <= 30'b000000010000000000100010110000
                ;mem[6526] <= 30'b000000010000000000100011010000
                ;mem[6527] <= 30'b000000010000000000100011100000
                ;mem[6528] <= 30'b000000010000000000100011110000
                ;mem[6529] <= 30'b000000010000000000101010010000
                ;mem[6530] <= 30'b000000010000000000101010100000
                ;mem[6531] <= 30'b000000010000000000110001010000
                ;mem[6532] <= 30'b000000010000000000110001100000
                ;mem[6533] <= 30'b000000010000000000110001110000
                ;mem[6534] <= 30'b000000010000000000111000010000
                ;mem[6535] <= 30'b000000010000000000111000100000
                ;mem[6536] <= 30'b000000010000000000111111010000
                ;mem[6537] <= 30'b000000010000000000111111100000
                ;mem[6538] <= 30'b000000000000000001000101010000
                ;mem[6539] <= 30'b000000000000000001000101100000
                ;mem[6540] <= 30'b000000000000000001000101110000
                ;mem[6541] <= 30'b000000000000000001001100010000
                ;mem[6542] <= 30'b000000000000000001001100100000
                ;mem[6543] <= 30'b000000000000000001010011010000
                ;mem[6544] <= 30'b000000000000000001010011100000
                ;mem[6545] <= 30'b000000000000000001011010010000
                ;mem[6546] <= 30'b000000000000000001011010100000
                ;mem[6547] <= 30'b000000000000000001100001010000
                ;mem[6548] <= 30'b000000000000000001100001100000
                ;mem[6549] <= 30'b000000000000000001101000100000
                ;mem[6550] <= 30'b000000000000000000011001010000
                ;mem[6551] <= 30'b000000000000000000011001100000
                ;mem[6552] <= 30'b000000000000000000100000000000
                ;mem[6553] <= 30'b000000000000000000100000010000
                ;mem[6554] <= 30'b000000000000000000100000100000
                ;mem[6555] <= 30'b000000000000000000100111000000
                ;mem[6556] <= 30'b000000000000000000100111010000
                ;mem[6557] <= 30'b000000000000000000100111100000
                ;mem[6558] <= 30'b000000000000000000101101110000
                ;mem[6559] <= 30'b000000000000000000101110000000
                ;mem[6560] <= 30'b000000000000000000101110010000
                ;mem[6561] <= 30'b000000000000000000110100100000
                ;mem[6562] <= 30'b000000000000000000110100110000
                ;mem[6563] <= 30'b000000000000000000110101000000
                ;mem[6564] <= 30'b000000000000000000111011100000
                ;mem[6565] <= 30'b000000000000000000111011110000
                ;mem[6566] <= 30'b000000001000000000000001110000
                ;mem[6567] <= 30'b000000001000000000000010000000
                ;mem[6568] <= 30'b000000001000000000000010010000
                ;mem[6569] <= 30'b000000001000000000001000100000
                ;mem[6570] <= 30'b000000001000000000001000110000
                ;mem[6571] <= 30'b000000001000000000001001000000
                ;mem[6572] <= 30'b000000001000000000001111100000
                ;mem[6573] <= 30'b000000001000000000001111110000
                ;mem[6574] <= 30'b000000001000000000010110010000
                ;mem[6575] <= 30'b000000001000000000010110100000
                ;mem[6576] <= 30'b000000001000000000011101010000
                ;mem[6577] <= 30'b000000001000000000011101100000
                ;mem[6578] <= 30'b000000001000000000100011110000
                ;mem[6579] <= 30'b000000001000000000100100000000
                ;mem[6580] <= 30'b000000001000000000100100010000
                ;mem[6581] <= 30'b000000001000000000101010110000
                ;mem[6582] <= 30'b000000001000000000101011000000
                ;mem[6583] <= 30'b000000001000000000110001100000
                ;mem[6584] <= 30'b000000001000000000110001110000
                ;mem[6585] <= 30'b000000001000000000110010000000
                ;mem[6586] <= 30'b000000001000000000111000100000
                ;mem[6587] <= 30'b000000001000000000111000110000
                ;mem[6588] <= 30'b000000001000000000111001110000
                ;mem[6589] <= 30'b000000001000000000111010000000
                ;mem[6590] <= 30'b000000001000000000111010010000
                ;mem[6591] <= 30'b000000001000000000111010100000
                ;mem[6592] <= 30'b000000001000000000111111100000
                ;mem[6593] <= 30'b000000001000000000111111110000
                ;mem[6594] <= 30'b000000010000000000000101100000
                ;mem[6595] <= 30'b000000010000000000000101110000
                ;mem[6596] <= 30'b000000010000000000000110000000
                ;mem[6597] <= 30'b000000010000000000001100100000
                ;mem[6598] <= 30'b000000010000000000001100110000
                ;mem[6599] <= 30'b000000010000000000001101110000
                ;mem[6600] <= 30'b000000010000000000001110000000
                ;mem[6601] <= 30'b000000010000000000001110010000
                ;mem[6602] <= 30'b000000010000000000001110100000
                ;mem[6603] <= 30'b000000010000000000010011100000
                ;mem[6604] <= 30'b000000010000000000010011110000
                ;mem[6605] <= 30'b000000010000000000010100100000
                ;mem[6606] <= 30'b000000010000000000010100110000
                ;mem[6607] <= 30'b000000010000000000010101000000
                ;mem[6608] <= 30'b000000010000000000010101010000
                ;mem[6609] <= 30'b000000010000000000010101100000
                ;mem[6610] <= 30'b000000010000000000010101110000
                ;mem[6611] <= 30'b000000010000000000011010010000
                ;mem[6612] <= 30'b000000010000000000011010100000
                ;mem[6613] <= 30'b000000010000000000011010110000
                ;mem[6614] <= 30'b000000010000000000011100010000
                ;mem[6615] <= 30'b000000010000000000011100100000
                ;mem[6616] <= 30'b000000010000000000011100110000
                ;mem[6617] <= 30'b000000010000000000100001010000
                ;mem[6618] <= 30'b000000010000000000100001100000
                ;mem[6619] <= 30'b000000010000000000100011010000
                ;mem[6620] <= 30'b000000010000000000100011100000
                ;mem[6621] <= 30'b000000010000000000100011110000
                ;mem[6622] <= 30'b000000010000000000101000010000
                ;mem[6623] <= 30'b000000010000000000101000100000
                ;mem[6624] <= 30'b000000010000000000101000110000
                ;mem[6625] <= 30'b000000010000000000101010010000
                ;mem[6626] <= 30'b000000010000000000101010100000
                ;mem[6627] <= 30'b000000010000000000101010110000
                ;mem[6628] <= 30'b000000010000000000101111010000
                ;mem[6629] <= 30'b000000010000000000101111100000
                ;mem[6630] <= 30'b000000010000000000101111110000
                ;mem[6631] <= 30'b000000010000000000110001010000
                ;mem[6632] <= 30'b000000010000000000110001100000
                ;mem[6633] <= 30'b000000010000000000110110010000
                ;mem[6634] <= 30'b000000010000000000110110100000
                ;mem[6635] <= 30'b000000010000000000110110110000
                ;mem[6636] <= 30'b000000010000000000110111000000
                ;mem[6637] <= 30'b000000010000000000110111010000
                ;mem[6638] <= 30'b000000010000000000110111110000
                ;mem[6639] <= 30'b000000010000000000111000000000
                ;mem[6640] <= 30'b000000010000000000111000010000
                ;mem[6641] <= 30'b000000010000000000111000100000
                ;mem[6642] <= 30'b000000010000000000111101110000
                ;mem[6643] <= 30'b000000010000000000111110000000
                ;mem[6644] <= 30'b000000010000000000111110010000
                ;mem[6645] <= 30'b000000010000000000111110100000
                ;mem[6646] <= 30'b000000010000000000111110110000
                ;mem[6647] <= 30'b000000010000000000111111000000
                ;mem[6648] <= 30'b000000010000000000111111010000
                ;mem[6649] <= 30'b000000000000000001000011010000
                ;mem[6650] <= 30'b000000000000000001000011100000
                ;mem[6651] <= 30'b000000000000000001000011110000
                ;mem[6652] <= 30'b000000000000000001000101010000
                ;mem[6653] <= 30'b000000000000000001000101100000
                ;mem[6654] <= 30'b000000000000000001001010010000
                ;mem[6655] <= 30'b000000000000000001001010100000
                ;mem[6656] <= 30'b000000000000000001001010110000
                ;mem[6657] <= 30'b000000000000000001001011000000
                ;mem[6658] <= 30'b000000000000000001001011010000
                ;mem[6659] <= 30'b000000000000000001001011110000
                ;mem[6660] <= 30'b000000000000000001001100000000
                ;mem[6661] <= 30'b000000000000000001001100010000
                ;mem[6662] <= 30'b000000000000000001001100100000
                ;mem[6663] <= 30'b000000000000000001010001110000
                ;mem[6664] <= 30'b000000000000000001010010000000
                ;mem[6665] <= 30'b000000000000000001010010010000
                ;mem[6666] <= 30'b000000000000000001010010100000
                ;mem[6667] <= 30'b000000000000000001010010110000
                ;mem[6668] <= 30'b000000000000000001010011000000
                ;mem[6669] <= 30'b000000000000000001010011010000
                ;mem[6670] <= 30'b000000000000000001011001010000
                ;mem[6671] <= 30'b000000000000000001011001100000
                ;mem[6672] <= 30'b000000000000000001011001110000
                ;mem[6673] <= 30'b000000000000000000101011110000
                ;mem[6674] <= 30'b000000000000000000101100000000
                ;mem[6675] <= 30'b000000000000000000101100010000
                ;mem[6676] <= 30'b000000000000000000101100100000
                ;mem[6677] <= 30'b000000000000000000101100110000
                ;mem[6678] <= 30'b000000000000000000101101000000
                ;mem[6679] <= 30'b000000000000000000101101010000
                ;mem[6680] <= 30'b000000000000000000101101100000
                ;mem[6681] <= 30'b000000000000000000101101110000
                ;mem[6682] <= 30'b000000000000000000110010000000
                ;mem[6683] <= 30'b000000000000000000110010010000
                ;mem[6684] <= 30'b000000000000000000110010100000
                ;mem[6685] <= 30'b000000000000000000110010110000
                ;mem[6686] <= 30'b000000000000000000110011000000
                ;mem[6687] <= 30'b000000000000000000110011010000
                ;mem[6688] <= 30'b000000000000000000110011100000
                ;mem[6689] <= 30'b000000000000000000110011110000
                ;mem[6690] <= 30'b000000000000000000110100000000
                ;mem[6691] <= 30'b000000000000000000110100010000
                ;mem[6692] <= 30'b000000000000000000110100100000
                ;mem[6693] <= 30'b000000000000000000110100110000
                ;mem[6694] <= 30'b000000000000000000110101000000
                ;mem[6695] <= 30'b000000000000000000110101010000
                ;mem[6696] <= 30'b000000000000000000111001000000
                ;mem[6697] <= 30'b000000000000000000111001010000
                ;mem[6698] <= 30'b000000000000000000111001100000
                ;mem[6699] <= 30'b000000000000000000111001110000
                ;mem[6700] <= 30'b000000000000000000111010000000
                ;mem[6701] <= 30'b000000000000000000111010010000
                ;mem[6702] <= 30'b000000000000000000111010100000
                ;mem[6703] <= 30'b000000000000000000111010110000
                ;mem[6704] <= 30'b000000000000000000111011000000
                ;mem[6705] <= 30'b000000000000000000111011010000
                ;mem[6706] <= 30'b000000000000000000111011100000
                ;mem[6707] <= 30'b000000000000000000111011110000
                ;mem[6708] <= 30'b000000000000000000111100000000
                ;mem[6709] <= 30'b000000000000000000111100010000
                ;mem[6710] <= 30'b000000000000000000111100100000
                ;mem[6711] <= 30'b000000001000000000000000000000
                ;mem[6712] <= 30'b000000001000000000000000010000
                ;mem[6713] <= 30'b000000001000000000000000100000
                ;mem[6714] <= 30'b000000001000000000000000110000
                ;mem[6715] <= 30'b000000001000000000000001000000
                ;mem[6716] <= 30'b000000001000000000000001010000
                ;mem[6717] <= 30'b000000001000000000000001100000
                ;mem[6718] <= 30'b000000001000000000000001110000
                ;mem[6719] <= 30'b000000001000000000000110000000
                ;mem[6720] <= 30'b000000001000000000000110010000
                ;mem[6721] <= 30'b000000001000000000000110100000
                ;mem[6722] <= 30'b000000001000000000000110110000
                ;mem[6723] <= 30'b000000001000000000000111000000
                ;mem[6724] <= 30'b000000001000000000000111010000
                ;mem[6725] <= 30'b000000001000000000000111100000
                ;mem[6726] <= 30'b000000001000000000000111110000
                ;mem[6727] <= 30'b000000001000000000001000000000
                ;mem[6728] <= 30'b000000001000000000001000010000
                ;mem[6729] <= 30'b000000001000000000001000100000
                ;mem[6730] <= 30'b000000001000000000001000110000
                ;mem[6731] <= 30'b000000001000000000001001000000
                ;mem[6732] <= 30'b000000001000000000001001010000
                ;mem[6733] <= 30'b000000001000000000001101000000
                ;mem[6734] <= 30'b000000001000000000001101010000
                ;mem[6735] <= 30'b000000001000000000001101100000
                ;mem[6736] <= 30'b000000001000000000001101110000
                ;mem[6737] <= 30'b000000001000000000001110000000
                ;mem[6738] <= 30'b000000001000000000001110010000
                ;mem[6739] <= 30'b000000001000000000001110100000
                ;mem[6740] <= 30'b000000001000000000001110110000
                ;mem[6741] <= 30'b000000001000000000001111000000
                ;mem[6742] <= 30'b000000001000000000001111010000
                ;mem[6743] <= 30'b000000001000000000001111100000
                ;mem[6744] <= 30'b000000001000000000001111110000
                ;mem[6745] <= 30'b000000001000000000010000000000
                ;mem[6746] <= 30'b000000001000000000010000010000
                ;mem[6747] <= 30'b000000001000000000010000100000
                ;mem[6748] <= 30'b000000001000000000010100010000
                ;mem[6749] <= 30'b000000001000000000010100100000
                ;mem[6750] <= 30'b000000001000000000010100110000
                ;mem[6751] <= 30'b000000001000000000010101000000
                ;mem[6752] <= 30'b000000001000000000010101010000
                ;mem[6753] <= 30'b000000001000000000010110110000
                ;mem[6754] <= 30'b000000001000000000010111000000
                ;mem[6755] <= 30'b000000001000000000010111010000
                ;mem[6756] <= 30'b000000001000000000010111100000
                ;mem[6757] <= 30'b000000001000000000011101110000
                ;mem[6758] <= 30'b000000001000000000011110000000
                ;mem[6759] <= 30'b000000001000000000011110010000
                ;mem[6760] <= 30'b000000001000000000011110100000
                ;mem[6761] <= 30'b000000001000000000100100010000
                ;mem[6762] <= 30'b000000001000000000100100100000
                ;mem[6763] <= 30'b000000001000000000100100110000
                ;mem[6764] <= 30'b000000001000000000100101000000
                ;mem[6765] <= 30'b000000001000000000100101010000
                ;mem[6766] <= 30'b000000001000000000101010110000
                ;mem[6767] <= 30'b000000001000000000101011000000
                ;mem[6768] <= 30'b000000001000000000101011010000
                ;mem[6769] <= 30'b000000001000000000101011100000
                ;mem[6770] <= 30'b000000001000000000101011110000
                ;mem[6771] <= 30'b000000001000000000101100000000
                ;mem[6772] <= 30'b000000001000000000101100010000
                ;mem[6773] <= 30'b000000001000000000110001000000
                ;mem[6774] <= 30'b000000001000000000110001010000
                ;mem[6775] <= 30'b000000001000000000110001100000
                ;mem[6776] <= 30'b000000001000000000110001110000
                ;mem[6777] <= 30'b000000001000000000110010000000
                ;mem[6778] <= 30'b000000001000000000110010010000
                ;mem[6779] <= 30'b000000001000000000110010100000
                ;mem[6780] <= 30'b000000001000000000110010110000
                ;mem[6781] <= 30'b000000001000000000110011000000
                ;mem[6782] <= 30'b000000001000000000110011010000
                ;mem[6783] <= 30'b000000001000000000110011100000
                ;mem[6784] <= 30'b000000001000000000110011110000
                ;mem[6785] <= 30'b000000001000000000111000000000
                ;mem[6786] <= 30'b000000001000000000111000010000
                ;mem[6787] <= 30'b000000001000000000111000100000
                ;mem[6788] <= 30'b000000001000000000111000110000
                ;mem[6789] <= 30'b000000001000000000111001000000
                ;mem[6790] <= 30'b000000001000000000111001010000
                ;mem[6791] <= 30'b000000001000000000111001100000
                ;mem[6792] <= 30'b000000001000000000111001110000
                ;mem[6793] <= 30'b000000001000000000111010000000
                ;mem[6794] <= 30'b000000001000000000111010010000
                ;mem[6795] <= 30'b000000001000000000111010100000
                ;mem[6796] <= 30'b000000001000000000111010110000
                ;mem[6797] <= 30'b000000001000000000111011000000
                ;mem[6798] <= 30'b000000001000000000111011010000
                ;mem[6799] <= 30'b000000001000000000111011100000
                ;mem[6800] <= 30'b000000001000000000111111000000
                ;mem[6801] <= 30'b000000001000000000111111010000
                ;mem[6802] <= 30'b000000001000000000111111100000
                ;mem[6803] <= 30'b000000001000000000111111110000
                ;mem[6804] <= 30'b000000010000000000000000000000
                ;mem[6805] <= 30'b000000010000000000000000010000
                ;mem[6806] <= 30'b000000010000000000000101000000
                ;mem[6807] <= 30'b000000010000000000000101010000
                ;mem[6808] <= 30'b000000010000000000000101100000
                ;mem[6809] <= 30'b000000010000000000000101110000
                ;mem[6810] <= 30'b000000010000000000000110000000
                ;mem[6811] <= 30'b000000010000000000000110010000
                ;mem[6812] <= 30'b000000010000000000000110100000
                ;mem[6813] <= 30'b000000010000000000000110110000
                ;mem[6814] <= 30'b000000010000000000000111000000
                ;mem[6815] <= 30'b000000010000000000000111010000
                ;mem[6816] <= 30'b000000010000000000000111100000
                ;mem[6817] <= 30'b000000010000000000000111110000
                ;mem[6818] <= 30'b000000010000000000001100000000
                ;mem[6819] <= 30'b000000010000000000001100010000
                ;mem[6820] <= 30'b000000010000000000001100100000
                ;mem[6821] <= 30'b000000010000000000001100110000
                ;mem[6822] <= 30'b000000010000000000001101000000
                ;mem[6823] <= 30'b000000010000000000001101010000
                ;mem[6824] <= 30'b000000010000000000001101100000
                ;mem[6825] <= 30'b000000010000000000001101110000
                ;mem[6826] <= 30'b000000010000000000001110000000
                ;mem[6827] <= 30'b000000010000000000001110010000
                ;mem[6828] <= 30'b000000010000000000001110100000
                ;mem[6829] <= 30'b000000010000000000001110110000
                ;mem[6830] <= 30'b000000010000000000001111000000
                ;mem[6831] <= 30'b000000010000000000001111010000
                ;mem[6832] <= 30'b000000010000000000001111100000
                ;mem[6833] <= 30'b000000010000000000010011000000
                ;mem[6834] <= 30'b000000010000000000010011010000
                ;mem[6835] <= 30'b000000010000000000010011100000
                ;mem[6836] <= 30'b000000010000000000010011110000
                ;mem[6837] <= 30'b000000010000000000010101100000
                ;mem[6838] <= 30'b000000010000000000010101110000
                ;mem[6839] <= 30'b000000010000000000010110000000
                ;mem[6840] <= 30'b000000010000000000010110010000
                ;mem[6841] <= 30'b000000010000000000010110100000
                ;mem[6842] <= 30'b000000010000000000011101000000
                ;mem[6843] <= 30'b000000010000000000011101010000
                ;mem[6844] <= 30'b000000010000000000011101100000
                ;mem[6845] <= 30'b000000010000000000011101110000
                ;mem[6846] <= 30'b000000010000000000100100010000
                ;mem[6847] <= 30'b000000010000000000100100100000
                ;mem[6848] <= 30'b000000010000000000100100110000
                ;mem[6849] <= 30'b000000010000000000101011010000
                ;mem[6850] <= 30'b000000010000000000101011100000
                ;mem[6851] <= 30'b000000010000000000101011110000
                ;mem[6852] <= 30'b000000010000000000101111010000
                ;mem[6853] <= 30'b000000010000000000101111100000
                ;mem[6854] <= 30'b000000010000000000110010000000
                ;mem[6855] <= 30'b000000010000000000110010010000
                ;mem[6856] <= 30'b000000010000000000110010100000
                ;mem[6857] <= 30'b000000010000000000110110010000
                ;mem[6858] <= 30'b000000010000000000110110100000
                ;mem[6859] <= 30'b000000010000000000110110110000
                ;mem[6860] <= 30'b000000010000000000110111000000
                ;mem[6861] <= 30'b000000010000000000110111010000
                ;mem[6862] <= 30'b000000010000000000111000000000
                ;mem[6863] <= 30'b000000010000000000111000010000
                ;mem[6864] <= 30'b000000010000000000111000100000
                ;mem[6865] <= 30'b000000010000000000111000110000
                ;mem[6866] <= 30'b000000010000000000111001000000
                ;mem[6867] <= 30'b000000010000000000111001010000
                ;mem[6868] <= 30'b000000010000000000111001100000
                ;mem[6869] <= 30'b000000010000000000111101010000
                ;mem[6870] <= 30'b000000010000000000111101100000
                ;mem[6871] <= 30'b000000010000000000111101110000
                ;mem[6872] <= 30'b000000010000000000111110000000
                ;mem[6873] <= 30'b000000010000000000111110010000
                ;mem[6874] <= 30'b000000010000000000111110100000
                ;mem[6875] <= 30'b000000010000000000111110110000
                ;mem[6876] <= 30'b000000010000000000111111000000
                ;mem[6877] <= 30'b000000010000000000111111010000
                ;mem[6878] <= 30'b000000010000000000111111100000
                ;mem[6879] <= 30'b000000010000000000111111110000
                ;mem[6880] <= 30'b000000000000000001000011010000
                ;mem[6881] <= 30'b000000000000000001000011100000
                ;mem[6882] <= 30'b000000000000000001000110000000
                ;mem[6883] <= 30'b000000000000000001000110010000
                ;mem[6884] <= 30'b000000000000000001000110100000
                ;mem[6885] <= 30'b000000000000000001001010010000
                ;mem[6886] <= 30'b000000000000000001001010100000
                ;mem[6887] <= 30'b000000000000000001001010110000
                ;mem[6888] <= 30'b000000000000000001001011000000
                ;mem[6889] <= 30'b000000000000000001001011010000
                ;mem[6890] <= 30'b000000000000000001001100000000
                ;mem[6891] <= 30'b000000000000000001001100010000
                ;mem[6892] <= 30'b000000000000000001001100100000
                ;mem[6893] <= 30'b000000000000000001001100110000
                ;mem[6894] <= 30'b000000000000000001001101000000
                ;mem[6895] <= 30'b000000000000000001001101010000
                ;mem[6896] <= 30'b000000000000000001001101100000
                ;mem[6897] <= 30'b000000000000000001010001010000
                ;mem[6898] <= 30'b000000000000000001010001100000
                ;mem[6899] <= 30'b000000000000000001010001110000
                ;mem[6900] <= 30'b000000000000000001010010000000
                ;mem[6901] <= 30'b000000000000000001010010010000
                ;mem[6902] <= 30'b000000000000000001010010100000
                ;mem[6903] <= 30'b000000000000000001010010110000
                ;mem[6904] <= 30'b000000000000000001010011000000
                ;mem[6905] <= 30'b000000000000000001010011010000
                ;mem[6906] <= 30'b000000000000000001010011100000
                ;mem[6907] <= 30'b000000000000000001010011110000
                ;mem[6908] <= 30'b000000000000000001010100000000
                ;mem[6909] <= 30'b000000000000000001010100010000
                ;mem[6910] <= 30'b000000000000000001011000110000
                ;mem[6911] <= 30'b000000000000000001011001000000
                ;mem[6912] <= 30'b000000000000000001011001010000
                ;mem[6913] <= 30'b000000000000000001011001100000
                ;mem[6914] <= 30'b000000000000000001011001110000
                ;mem[6915] <= 30'b000000000000000001011010000000
                ;mem[6916] <= 30'b000000000000000001011010010000
                ;mem[6917] <= 30'b000000000000000001011010100000
                ;mem[6918] <= 30'b000000000000000001011010110000
                ;mem[6919] <= 30'b000000000000000001011011000000
                ;mem[6920] <= 30'b000000000000000000101111010000
                ;mem[6921] <= 30'b000000000000000000101111100000
                ;mem[6922] <= 30'b000000000000000000101111110000
                ;mem[6923] <= 30'b000000000000000000110000000000
                ;mem[6924] <= 30'b000000000000000000110101100000
                ;mem[6925] <= 30'b000000000000000000110101110000
                ;mem[6926] <= 30'b000000000000000000110110000000
                ;mem[6927] <= 30'b000000000000000000110110010000
                ;mem[6928] <= 30'b000000000000000000110110100000
                ;mem[6929] <= 30'b000000000000000000111011000000
                ;mem[6930] <= 30'b000000000000000000111011010000
                ;mem[6931] <= 30'b000000000000000000111011100000
                ;mem[6932] <= 30'b000000000000000000111011110000
                ;mem[6933] <= 30'b000000000000000000111100000000
                ;mem[6934] <= 30'b000000000000000000111100010000
                ;mem[6935] <= 30'b000000000000000000111100100000
                ;mem[6936] <= 30'b000000000000000000111100110000
                ;mem[6937] <= 30'b000000001000000000000011010000
                ;mem[6938] <= 30'b000000001000000000000011100000
                ;mem[6939] <= 30'b000000001000000000000011110000
                ;mem[6940] <= 30'b000000001000000000000100000000
                ;mem[6941] <= 30'b000000001000000000001001100000
                ;mem[6942] <= 30'b000000001000000000001001110000
                ;mem[6943] <= 30'b000000001000000000001010000000
                ;mem[6944] <= 30'b000000001000000000001010010000
                ;mem[6945] <= 30'b000000001000000000001010100000
                ;mem[6946] <= 30'b000000001000000000001111000000
                ;mem[6947] <= 30'b000000001000000000001111010000
                ;mem[6948] <= 30'b000000001000000000001111100000
                ;mem[6949] <= 30'b000000001000000000001111110000
                ;mem[6950] <= 30'b000000001000000000010000000000
                ;mem[6951] <= 30'b000000001000000000010000010000
                ;mem[6952] <= 30'b000000001000000000010000100000
                ;mem[6953] <= 30'b000000001000000000010000110000
                ;mem[6954] <= 30'b000000001000000000010101110000
                ;mem[6955] <= 30'b000000001000000000010110000000
                ;mem[6956] <= 30'b000000001000000000010110010000
                ;mem[6957] <= 30'b000000001000000000010110100000
                ;mem[6958] <= 30'b000000001000000000010110110000
                ;mem[6959] <= 30'b000000001000000000010111000000
                ;mem[6960] <= 30'b000000001000000000011100100000
                ;mem[6961] <= 30'b000000001000000000011100110000
                ;mem[6962] <= 30'b000000001000000000011101000000
                ;mem[6963] <= 30'b000000001000000000011101010000
                ;mem[6964] <= 30'b000000001000000000011101100000
                ;mem[6965] <= 30'b000000001000000000100011010000
                ;mem[6966] <= 30'b000000001000000000100011100000
                ;mem[6967] <= 30'b000000001000000000100011110000
                ;mem[6968] <= 30'b000000001000000000100100000000
                ;mem[6969] <= 30'b000000001000000000101010010000
                ;mem[6970] <= 30'b000000001000000000101010100000
                ;mem[6971] <= 30'b000000001000000000101010110000
                ;mem[6972] <= 30'b000000001000000000110001000000
                ;mem[6973] <= 30'b000000001000000000110001010000
                ;mem[6974] <= 30'b000000001000000000110001100000
                ;mem[6975] <= 30'b000000001000000000111000000000
                ;mem[6976] <= 30'b000000001000000000111000010000
                ;mem[6977] <= 30'b000000001000000000111001010000
                ;mem[6978] <= 30'b000000001000000000111001100000
                ;mem[6979] <= 30'b000000001000000000111001110000
                ;mem[6980] <= 30'b000000001000000000111111000000
                ;mem[6981] <= 30'b000000001000000000111111010000
                ;mem[6982] <= 30'b000000001000000000111111100000
                ;mem[6983] <= 30'b000000001000000000111111110000
                ;mem[6984] <= 30'b000000010000000000000101000000
                ;mem[6985] <= 30'b000000010000000000000101010000
                ;mem[6986] <= 30'b000000010000000000000101100000
                ;mem[6987] <= 30'b000000010000000000001100000000
                ;mem[6988] <= 30'b000000010000000000001100010000
                ;mem[6989] <= 30'b000000010000000000001101010000
                ;mem[6990] <= 30'b000000010000000000001101100000
                ;mem[6991] <= 30'b000000010000000000001101110000
                ;mem[6992] <= 30'b000000010000000000010011000000
                ;mem[6993] <= 30'b000000010000000000010011010000
                ;mem[6994] <= 30'b000000010000000000010011100000
                ;mem[6995] <= 30'b000000010000000000010011110000
                ;mem[6996] <= 30'b000000010000000000010100000000
                ;mem[6997] <= 30'b000000010000000000010100010000
                ;mem[6998] <= 30'b000000010000000000010100100000
                ;mem[6999] <= 30'b000000010000000000010100110000
                ;mem[7000] <= 30'b000000010000000000010101000000
                ;mem[7001] <= 30'b000000010000000000010101010000
                ;mem[7002] <= 30'b000000010000000000011001110000
                ;mem[7003] <= 30'b000000010000000000011010000000
                ;mem[7004] <= 30'b000000010000000000011010010000
                ;mem[7005] <= 30'b000000010000000000011010100000
                ;mem[7006] <= 30'b000000010000000000011010110000
                ;mem[7007] <= 30'b000000010000000000011100000000
                ;mem[7008] <= 30'b000000010000000000011100010000
                ;mem[7009] <= 30'b000000010000000000011100100000
                ;mem[7010] <= 30'b000000010000000000100001000000
                ;mem[7011] <= 30'b000000010000000000100011010000
                ;mem[7012] <= 30'b000000010000000000100011100000
                ;mem[7013] <= 30'b000000010000000000100011110000
                ;mem[7014] <= 30'b000000010000000000101010100000
                ;mem[7015] <= 30'b000000010000000000101010110000
                ;mem[7016] <= 30'b000000010000000000110001010000
                ;mem[7017] <= 30'b000000010000000000110001100000
                ;mem[7018] <= 30'b000000010000000000110001110000
                ;mem[7019] <= 30'b000000010000000000111000000000
                ;mem[7020] <= 30'b000000010000000000111000010000
                ;mem[7021] <= 30'b000000010000000000111000100000
                ;mem[7022] <= 30'b000000010000000000111110100000
                ;mem[7023] <= 30'b000000010000000000111110110000
                ;mem[7024] <= 30'b000000010000000000111111000000
                ;mem[7025] <= 30'b000000010000000000111111010000
                ;mem[7026] <= 30'b000000000000000001000101010000
                ;mem[7027] <= 30'b000000000000000001000101100000
                ;mem[7028] <= 30'b000000000000000001000101110000
                ;mem[7029] <= 30'b000000000000000001001100000000
                ;mem[7030] <= 30'b000000000000000001001100010000
                ;mem[7031] <= 30'b000000000000000001001100100000
                ;mem[7032] <= 30'b000000000000000001010010100000
                ;mem[7033] <= 30'b000000000000000001010010110000
                ;mem[7034] <= 30'b000000000000000001010011000000
                ;mem[7035] <= 30'b000000000000000001010011010000
                ;mem[7036] <= 30'b000000000000000001011000110000
                ;mem[7037] <= 30'b000000000000000001011001000000
                ;mem[7038] <= 30'b000000000000000001011001010000
                ;mem[7039] <= 30'b000000000000000001011001100000
                ;mem[7040] <= 30'b000000000000000001011001110000
                ;mem[7041] <= 30'b000000000000000001011010000000
                ;mem[7042] <= 30'b000000000000000001011110100000
                ;mem[7043] <= 30'b000000000000000001011110110000
                ;mem[7044] <= 30'b000000000000000001011111000000
                ;mem[7045] <= 30'b000000000000000001011111010000
                ;mem[7046] <= 30'b000000000000000001011111100000
                ;mem[7047] <= 30'b000000000000000001011111110000
                ;mem[7048] <= 30'b000000000000000001100000000000
                ;mem[7049] <= 30'b000000000000000001100000010000
                ;mem[7050] <= 30'b000000000000000000011111110000
                ;mem[7051] <= 30'b000000000000000000100000000000
                ;mem[7052] <= 30'b000000000000000000100000010000
                ;mem[7053] <= 30'b000000000000000000100110100000
                ;mem[7054] <= 30'b000000000000000000100110110000
                ;mem[7055] <= 30'b000000000000000000101100010000
                ;mem[7056] <= 30'b000000000000000000101100100000
                ;mem[7057] <= 30'b000000000000000000101100110000
                ;mem[7058] <= 30'b000000000000000000101101000000
                ;mem[7059] <= 30'b000000000000000000101101010000
                ;mem[7060] <= 30'b000000000000000000110011000000
                ;mem[7061] <= 30'b000000000000000000110011010000
                ;mem[7062] <= 30'b000000000000000000110011100000
                ;mem[7063] <= 30'b000000000000000000110011110000
                ;mem[7064] <= 30'b000000000000000000111010000000
                ;mem[7065] <= 30'b000000001000000000000000010000
                ;mem[7066] <= 30'b000000001000000000000000100000
                ;mem[7067] <= 30'b000000001000000000000000110000
                ;mem[7068] <= 30'b000000001000000000000001000000
                ;mem[7069] <= 30'b000000001000000000000001010000
                ;mem[7070] <= 30'b000000001000000000000111000000
                ;mem[7071] <= 30'b000000001000000000000111010000
                ;mem[7072] <= 30'b000000001000000000000111100000
                ;mem[7073] <= 30'b000000001000000000000111110000
                ;mem[7074] <= 30'b000000001000000000001110000000
                ;mem[7075] <= 30'b000000001000000000010101000000
                ;mem[7076] <= 30'b000000001000000000011100000000
                ;mem[7077] <= 30'b000000001000000000100010110000
                ;mem[7078] <= 30'b000000001000000000100011000000
                ;mem[7079] <= 30'b000000001000000000101010000000
                ;mem[7080] <= 30'b000000001000000000101011000000
                ;mem[7081] <= 30'b000000001000000000101011010000
                ;mem[7082] <= 30'b000000001000000000101011100000
                ;mem[7083] <= 30'b000000001000000000101011110000
                ;mem[7084] <= 30'b000000001000000000101100000000
                ;mem[7085] <= 30'b000000001000000000101100010000
                ;mem[7086] <= 30'b000000001000000000101100100000
                ;mem[7087] <= 30'b000000001000000000110001000000
                ;mem[7088] <= 30'b000000001000000000110001010000
                ;mem[7089] <= 30'b000000001000000000110001100000
                ;mem[7090] <= 30'b000000001000000000110001110000
                ;mem[7091] <= 30'b000000001000000000110010000000
                ;mem[7092] <= 30'b000000001000000000110011100000
                ;mem[7093] <= 30'b000000001000000000110011110000
                ;mem[7094] <= 30'b000000001000000000111000000000
                ;mem[7095] <= 30'b000000001000000000111000010000
                ;mem[7096] <= 30'b000000001000000000111000100000
                ;mem[7097] <= 30'b000000001000000000111011000000
                ;mem[7098] <= 30'b000000010000000000000000000000
                ;mem[7099] <= 30'b000000010000000000000000010000
                ;mem[7100] <= 30'b000000010000000000000000100000
                ;mem[7101] <= 30'b000000010000000000000101000000
                ;mem[7102] <= 30'b000000010000000000000101010000
                ;mem[7103] <= 30'b000000010000000000000101100000
                ;mem[7104] <= 30'b000000010000000000000101110000
                ;mem[7105] <= 30'b000000010000000000000110000000
                ;mem[7106] <= 30'b000000010000000000000111100000
                ;mem[7107] <= 30'b000000010000000000000111110000
                ;mem[7108] <= 30'b000000010000000000001100000000
                ;mem[7109] <= 30'b000000010000000000001100010000
                ;mem[7110] <= 30'b000000010000000000001100100000
                ;mem[7111] <= 30'b000000010000000000001111000000
                ;mem[7112] <= 30'b000000010000000000010110000000
                ;mem[7113] <= 30'b000000010000000000010110010000
                ;mem[7114] <= 30'b000000010000000000011101010000
                ;mem[7115] <= 30'b000000010000000000100100010000
                ;mem[7116] <= 30'b000000010000000000101011010000
                ;mem[7117] <= 30'b000000010000000000110010000000
                ;mem[7118] <= 30'b000000010000000000110010010000
                ;mem[7119] <= 30'b000000010000000000111001000000
                ;mem[7120] <= 30'b000000010000000000111001010000
                ;mem[7121] <= 30'b000000010000000000111101010000
                ;mem[7122] <= 30'b000000010000000000111111100000
                ;mem[7123] <= 30'b000000010000000000111111110000
                ;mem[7124] <= 30'b000000000000000001000110000000
                ;mem[7125] <= 30'b000000000000000001000110010000
                ;mem[7126] <= 30'b000000000000000001001101000000
                ;mem[7127] <= 30'b000000000000000001001101010000
                ;mem[7128] <= 30'b000000000000000001010001010000
                ;mem[7129] <= 30'b000000000000000001010011100000
                ;mem[7130] <= 30'b000000000000000001010011110000
                ;mem[7131] <= 30'b000000000000000001010100000000
                ;mem[7132] <= 30'b000000000000000001011000100000
                ;mem[7133] <= 30'b000000000000000001011010000000
                ;mem[7134] <= 30'b000000000000000001011010010000
                ;mem[7135] <= 30'b000000000000000001011010100000
                ;mem[7136] <= 30'b000000000000000001011010110000
                ;mem[7137] <= 30'b000000000000000001011111100000
                ;mem[7138] <= 30'b000000000000000001011111110000
                ;mem[7139] <= 30'b000000000000000001100000000000
                ;mem[7140] <= 30'b000000000000000001100000010000
                ;mem[7141] <= 30'b000000000000000001100000100000
                ;mem[7142] <= 30'b000000000000000001100000110000
                ;mem[7143] <= 30'b000000000000000001100001000000
                ;mem[7144] <= 30'b000000000000000000010111100000
                ;mem[7145] <= 30'b000000000000000000010111110000
                ;mem[7146] <= 30'b000000000000000000011110010000
                ;mem[7147] <= 30'b000000000000000000011110100000
                ;mem[7148] <= 30'b000000000000000000011110110000
                ;mem[7149] <= 30'b000000000000000000100101000000
                ;mem[7150] <= 30'b000000000000000000100101010000
                ;mem[7151] <= 30'b000000000000000000100101100000
                ;mem[7152] <= 30'b000000000000000000100101110000
                ;mem[7153] <= 30'b000000000000000000101011110000
                ;mem[7154] <= 30'b000000000000000000101100000000
                ;mem[7155] <= 30'b000000000000000000101100010000
                ;mem[7156] <= 30'b000000000000000000101100100000
                ;mem[7157] <= 30'b000000000000000000110010110000
                ;mem[7158] <= 30'b000000000000000000110011000000
                ;mem[7159] <= 30'b000000000000000000110011010000
                ;mem[7160] <= 30'b000000000000000000111001100000
                ;mem[7161] <= 30'b000000000000000000111001110000
                ;mem[7162] <= 30'b000000000000000000111010000000
                ;mem[7163] <= 30'b000000000000000000111010010000
                ;mem[7164] <= 30'b000000001000000000000000000000
                ;mem[7165] <= 30'b000000001000000000000000010000
                ;mem[7166] <= 30'b000000001000000000000000100000
                ;mem[7167] <= 30'b000000001000000000000110110000
                ;mem[7168] <= 30'b000000001000000000000111000000
                ;mem[7169] <= 30'b000000001000000000000111010000
                ;mem[7170] <= 30'b000000001000000000001101100000
                ;mem[7171] <= 30'b000000001000000000001101110000
                ;mem[7172] <= 30'b000000001000000000001110000000
                ;mem[7173] <= 30'b000000001000000000001110010000
                ;mem[7174] <= 30'b000000001000000000010100100000
                ;mem[7175] <= 30'b000000001000000000010100110000
                ;mem[7176] <= 30'b000000001000000000010101000000
                ;mem[7177] <= 30'b000000001000000000011011100000
                ;mem[7178] <= 30'b000000001000000000011011110000
                ;mem[7179] <= 30'b000000001000000000011100000000
                ;mem[7180] <= 30'b000000001000000000100010100000
                ;mem[7181] <= 30'b000000001000000000100010110000
                ;mem[7182] <= 30'b000000001000000000100011000000
                ;mem[7183] <= 30'b000000001000000000100100110000
                ;mem[7184] <= 30'b000000001000000000100101000000
                ;mem[7185] <= 30'b000000001000000000100101010000
                ;mem[7186] <= 30'b000000001000000000100101100000
                ;mem[7187] <= 30'b000000001000000000100101110000
                ;mem[7188] <= 30'b000000001000000000100110000000
                ;mem[7189] <= 30'b000000001000000000100110010000
                ;mem[7190] <= 30'b000000001000000000100110100000
                ;mem[7191] <= 30'b000000001000000000101001100000
                ;mem[7192] <= 30'b000000001000000000101001110000
                ;mem[7193] <= 30'b000000001000000000101010000000
                ;mem[7194] <= 30'b000000001000000000101011100000
                ;mem[7195] <= 30'b000000001000000000101011110000
                ;mem[7196] <= 30'b000000001000000000101100000000
                ;mem[7197] <= 30'b000000001000000000101100010000
                ;mem[7198] <= 30'b000000001000000000101100100000
                ;mem[7199] <= 30'b000000001000000000101100110000
                ;mem[7200] <= 30'b000000001000000000101101000000
                ;mem[7201] <= 30'b000000001000000000101101010000
                ;mem[7202] <= 30'b000000001000000000101101100000
                ;mem[7203] <= 30'b000000001000000000101101110000
                ;mem[7204] <= 30'b000000001000000000101110000000
                ;mem[7205] <= 30'b000000001000000000110000100000
                ;mem[7206] <= 30'b000000001000000000110000110000
                ;mem[7207] <= 30'b000000001000000000110001000000
                ;mem[7208] <= 30'b000000001000000000110010010000
                ;mem[7209] <= 30'b000000001000000000110010100000
                ;mem[7210] <= 30'b000000001000000000110010110000
                ;mem[7211] <= 30'b000000001000000000110011000000
                ;mem[7212] <= 30'b000000001000000000110100110000
                ;mem[7213] <= 30'b000000001000000000110101000000
                ;mem[7214] <= 30'b000000001000000000110101010000
                ;mem[7215] <= 30'b000000001000000000110111100000
                ;mem[7216] <= 30'b000000001000000000110111110000
                ;mem[7217] <= 30'b000000001000000000111000000000
                ;mem[7218] <= 30'b000000001000000000111001010000
                ;mem[7219] <= 30'b000000001000000000111001100000
                ;mem[7220] <= 30'b000000001000000000111001110000
                ;mem[7221] <= 30'b000000001000000000111100000000
                ;mem[7222] <= 30'b000000001000000000111100010000
                ;mem[7223] <= 30'b000000001000000000111110100000
                ;mem[7224] <= 30'b000000001000000000111110110000
                ;mem[7225] <= 30'b000000001000000000111111000000
                ;mem[7226] <= 30'b000000010000000000000000000000
                ;mem[7227] <= 30'b000000010000000000000000010000
                ;mem[7228] <= 30'b000000010000000000000000100000
                ;mem[7229] <= 30'b000000010000000000000000110000
                ;mem[7230] <= 30'b000000010000000000000001000000
                ;mem[7231] <= 30'b000000010000000000000001010000
                ;mem[7232] <= 30'b000000010000000000000001100000
                ;mem[7233] <= 30'b000000010000000000000001110000
                ;mem[7234] <= 30'b000000010000000000000010000000
                ;mem[7235] <= 30'b000000010000000000000100100000
                ;mem[7236] <= 30'b000000010000000000000100110000
                ;mem[7237] <= 30'b000000010000000000000101000000
                ;mem[7238] <= 30'b000000010000000000000110010000
                ;mem[7239] <= 30'b000000010000000000000110100000
                ;mem[7240] <= 30'b000000010000000000000110110000
                ;mem[7241] <= 30'b000000010000000000000111000000
                ;mem[7242] <= 30'b000000010000000000001000110000
                ;mem[7243] <= 30'b000000010000000000001001000000
                ;mem[7244] <= 30'b000000010000000000001001010000
                ;mem[7245] <= 30'b000000010000000000001011100000
                ;mem[7246] <= 30'b000000010000000000001011110000
                ;mem[7247] <= 30'b000000010000000000001100000000
                ;mem[7248] <= 30'b000000010000000000001101010000
                ;mem[7249] <= 30'b000000010000000000001101100000
                ;mem[7250] <= 30'b000000010000000000001101110000
                ;mem[7251] <= 30'b000000010000000000010000000000
                ;mem[7252] <= 30'b000000010000000000010000010000
                ;mem[7253] <= 30'b000000010000000000010010100000
                ;mem[7254] <= 30'b000000010000000000010010110000
                ;mem[7255] <= 30'b000000010000000000010011000000
                ;mem[7256] <= 30'b000000010000000000010100010000
                ;mem[7257] <= 30'b000000010000000000010100100000
                ;mem[7258] <= 30'b000000010000000000010100110000
                ;mem[7259] <= 30'b000000010000000000010111000000
                ;mem[7260] <= 30'b000000010000000000010111010000
                ;mem[7261] <= 30'b000000010000000000011001100000
                ;mem[7262] <= 30'b000000010000000000011001110000
                ;mem[7263] <= 30'b000000010000000000011010000000
                ;mem[7264] <= 30'b000000010000000000011011010000
                ;mem[7265] <= 30'b000000010000000000011011100000
                ;mem[7266] <= 30'b000000010000000000011011110000
                ;mem[7267] <= 30'b000000010000000000011100000000
                ;mem[7268] <= 30'b000000010000000000011110000000
                ;mem[7269] <= 30'b000000010000000000100000110000
                ;mem[7270] <= 30'b000000010000000000100001000000
                ;mem[7271] <= 30'b000000010000000000100001010000
                ;mem[7272] <= 30'b000000010000000000100010110000
                ;mem[7273] <= 30'b000000010000000000100011000000
                ;mem[7274] <= 30'b000000010000000000100011010000
                ;mem[7275] <= 30'b000000010000000000100100110000
                ;mem[7276] <= 30'b000000010000000000100101000000
                ;mem[7277] <= 30'b000000010000000000100111110000
                ;mem[7278] <= 30'b000000010000000000101000000000
                ;mem[7279] <= 30'b000000010000000000101000010000
                ;mem[7280] <= 30'b000000010000000000101000100000
                ;mem[7281] <= 30'b000000010000000000101010000000
                ;mem[7282] <= 30'b000000010000000000101010010000
                ;mem[7283] <= 30'b000000010000000000101010100000
                ;mem[7284] <= 30'b000000010000000000101011110000
                ;mem[7285] <= 30'b000000010000000000101100000000
                ;mem[7286] <= 30'b000000010000000000101111000000
                ;mem[7287] <= 30'b000000010000000000101111010000
                ;mem[7288] <= 30'b000000010000000000101111100000
                ;mem[7289] <= 30'b000000010000000000101111110000
                ;mem[7290] <= 30'b000000010000000000110001010000
                ;mem[7291] <= 30'b000000010000000000110001100000
                ;mem[7292] <= 30'b000000010000000000110001110000
                ;mem[7293] <= 30'b000000010000000000110010000000
                ;mem[7294] <= 30'b000000010000000000110010100000
                ;mem[7295] <= 30'b000000010000000000110010110000
                ;mem[7296] <= 30'b000000010000000000110110010000
                ;mem[7297] <= 30'b000000010000000000110110100000
                ;mem[7298] <= 30'b000000010000000000110110110000
                ;mem[7299] <= 30'b000000010000000000110111000000
                ;mem[7300] <= 30'b000000010000000000110111010000
                ;mem[7301] <= 30'b000000010000000000111000110000
                ;mem[7302] <= 30'b000000010000000000111001000000
                ;mem[7303] <= 30'b000000010000000000111001010000
                ;mem[7304] <= 30'b000000010000000000111001100000
                ;mem[7305] <= 30'b000000010000000000111101100000
                ;mem[7306] <= 30'b000000010000000000111101110000
                ;mem[7307] <= 30'b000000010000000000111110000000
                ;mem[7308] <= 30'b000000010000000000111110010000
                ;mem[7309] <= 30'b000000010000000000111110100000
                ;mem[7310] <= 30'b000000010000000000111110110000
                ;mem[7311] <= 30'b000000010000000000111111000000
                ;mem[7312] <= 30'b000000010000000000111111010000
                ;mem[7313] <= 30'b000000010000000000111111100000
                ;mem[7314] <= 30'b000000010000000000111111110000
                ;mem[7315] <= 30'b000000000000000001000000000000
                ;mem[7316] <= 30'b000000000000000001000011000000
                ;mem[7317] <= 30'b000000000000000001000011010000
                ;mem[7318] <= 30'b000000000000000001000011100000
                ;mem[7319] <= 30'b000000000000000001000011110000
                ;mem[7320] <= 30'b000000000000000001000101010000
                ;mem[7321] <= 30'b000000000000000001000101100000
                ;mem[7322] <= 30'b000000000000000001000101110000
                ;mem[7323] <= 30'b000000000000000001000110000000
                ;mem[7324] <= 30'b000000000000000001000110100000
                ;mem[7325] <= 30'b000000000000000001000110110000
                ;mem[7326] <= 30'b000000000000000001001010010000
                ;mem[7327] <= 30'b000000000000000001001010100000
                ;mem[7328] <= 30'b000000000000000001001010110000
                ;mem[7329] <= 30'b000000000000000001001011000000
                ;mem[7330] <= 30'b000000000000000001001011010000
                ;mem[7331] <= 30'b000000000000000001001100110000
                ;mem[7332] <= 30'b000000000000000001001101000000
                ;mem[7333] <= 30'b000000000000000001001101010000
                ;mem[7334] <= 30'b000000000000000001001101100000
                ;mem[7335] <= 30'b000000000000000001010001100000
                ;mem[7336] <= 30'b000000000000000001010001110000
                ;mem[7337] <= 30'b000000000000000001010010000000
                ;mem[7338] <= 30'b000000000000000001010010010000
                ;mem[7339] <= 30'b000000000000000001010010100000
                ;mem[7340] <= 30'b000000000000000001010010110000
                ;mem[7341] <= 30'b000000000000000001010011000000
                ;mem[7342] <= 30'b000000000000000001010011010000
                ;mem[7343] <= 30'b000000000000000001010011100000
                ;mem[7344] <= 30'b000000000000000001010011110000
                ;mem[7345] <= 30'b000000000000000001010100000000
                ;mem[7346] <= 30'b000000000000000001011001010000
                ;mem[7347] <= 30'b000000000000000001011001100000
                ;mem[7348] <= 30'b000000000000000001011001110000
                ;mem[7349] <= 30'b000000000000000001011010000000
                ;mem[7350] <= 30'b000000000000000001011010010000
                ;mem[7351] <= 30'b000000000000000001011010100000
                ;mem[7352] <= 30'b000000000000000000100110110000
                ;mem[7353] <= 30'b000000000000000000100111000000
                ;mem[7354] <= 30'b000000000000000000100111010000
                ;mem[7355] <= 30'b000000000000000000101101000000
                ;mem[7356] <= 30'b000000000000000000101101010000
                ;mem[7357] <= 30'b000000000000000000101101100000
                ;mem[7358] <= 30'b000000000000000000101101110000
                ;mem[7359] <= 30'b000000000000000000101110000000
                ;mem[7360] <= 30'b000000000000000000101110010000
                ;mem[7361] <= 30'b000000000000000000110100000000
                ;mem[7362] <= 30'b000000000000000000110100010000
                ;mem[7363] <= 30'b000000000000000000110100100000
                ;mem[7364] <= 30'b000000000000000000110100110000
                ;mem[7365] <= 30'b000000000000000000110101010000
                ;mem[7366] <= 30'b000000000000000000110101100000
                ;mem[7367] <= 30'b000000000000000000110101110000
                ;mem[7368] <= 30'b000000000000000000111010110000
                ;mem[7369] <= 30'b000000000000000000111011000000
                ;mem[7370] <= 30'b000000000000000000111011010000
                ;mem[7371] <= 30'b000000000000000000111100010000
                ;mem[7372] <= 30'b000000000000000000111100100000
                ;mem[7373] <= 30'b000000000000000000111100110000
                ;mem[7374] <= 30'b000000001000000000000001000000
                ;mem[7375] <= 30'b000000001000000000000001010000
                ;mem[7376] <= 30'b000000001000000000000001100000
                ;mem[7377] <= 30'b000000001000000000000001110000
                ;mem[7378] <= 30'b000000001000000000000010000000
                ;mem[7379] <= 30'b000000001000000000000010010000
                ;mem[7380] <= 30'b000000001000000000001000000000
                ;mem[7381] <= 30'b000000001000000000001000010000
                ;mem[7382] <= 30'b000000001000000000001000100000
                ;mem[7383] <= 30'b000000001000000000001000110000
                ;mem[7384] <= 30'b000000001000000000001001010000
                ;mem[7385] <= 30'b000000001000000000001001100000
                ;mem[7386] <= 30'b000000001000000000001001110000
                ;mem[7387] <= 30'b000000001000000000001110110000
                ;mem[7388] <= 30'b000000001000000000001111000000
                ;mem[7389] <= 30'b000000001000000000001111010000
                ;mem[7390] <= 30'b000000001000000000010000010000
                ;mem[7391] <= 30'b000000001000000000010000100000
                ;mem[7392] <= 30'b000000001000000000010000110000
                ;mem[7393] <= 30'b000000001000000000010101100000
                ;mem[7394] <= 30'b000000001000000000010101110000
                ;mem[7395] <= 30'b000000001000000000010110000000
                ;mem[7396] <= 30'b000000001000000000010110010000
                ;mem[7397] <= 30'b000000001000000000010111100000
                ;mem[7398] <= 30'b000000001000000000010111110000
                ;mem[7399] <= 30'b000000001000000000011100100000
                ;mem[7400] <= 30'b000000001000000000011100110000
                ;mem[7401] <= 30'b000000001000000000011101000000
                ;mem[7402] <= 30'b000000001000000000011101010000
                ;mem[7403] <= 30'b000000001000000000011110100000
                ;mem[7404] <= 30'b000000001000000000011110110000
                ;mem[7405] <= 30'b000000001000000000011111000000
                ;mem[7406] <= 30'b000000001000000000100011100000
                ;mem[7407] <= 30'b000000001000000000100011110000
                ;mem[7408] <= 30'b000000001000000000100100000000
                ;mem[7409] <= 30'b000000001000000000100101110000
                ;mem[7410] <= 30'b000000001000000000100110000000
                ;mem[7411] <= 30'b000000001000000000101010100000
                ;mem[7412] <= 30'b000000001000000000101010110000
                ;mem[7413] <= 30'b000000001000000000101011000000
                ;mem[7414] <= 30'b000000001000000000101100110000
                ;mem[7415] <= 30'b000000001000000000101101000000
                ;mem[7416] <= 30'b000000001000000000110001100000
                ;mem[7417] <= 30'b000000001000000000110001110000
                ;mem[7418] <= 30'b000000001000000000110010000000
                ;mem[7419] <= 30'b000000001000000000110011110000
                ;mem[7420] <= 30'b000000001000000000110100000000
                ;mem[7421] <= 30'b000000001000000000111000010000
                ;mem[7422] <= 30'b000000001000000000111000100000
                ;mem[7423] <= 30'b000000001000000000111000110000
                ;mem[7424] <= 30'b000000001000000000111001000000
                ;mem[7425] <= 30'b000000001000000000111010110000
                ;mem[7426] <= 30'b000000001000000000111011000000
                ;mem[7427] <= 30'b000000001000000000111111010000
                ;mem[7428] <= 30'b000000001000000000111111100000
                ;mem[7429] <= 30'b000000001000000000111111110000
                ;mem[7430] <= 30'b000000010000000000000000110000
                ;mem[7431] <= 30'b000000010000000000000001000000
                ;mem[7432] <= 30'b000000010000000000000101100000
                ;mem[7433] <= 30'b000000010000000000000101110000
                ;mem[7434] <= 30'b000000010000000000000110000000
                ;mem[7435] <= 30'b000000010000000000000111110000
                ;mem[7436] <= 30'b000000010000000000001000000000
                ;mem[7437] <= 30'b000000010000000000001100010000
                ;mem[7438] <= 30'b000000010000000000001100100000
                ;mem[7439] <= 30'b000000010000000000001100110000
                ;mem[7440] <= 30'b000000010000000000001101000000
                ;mem[7441] <= 30'b000000010000000000001110110000
                ;mem[7442] <= 30'b000000010000000000001111000000
                ;mem[7443] <= 30'b000000010000000000010011010000
                ;mem[7444] <= 30'b000000010000000000010011100000
                ;mem[7445] <= 30'b000000010000000000010011110000
                ;mem[7446] <= 30'b000000010000000000010100000000
                ;mem[7447] <= 30'b000000010000000000010101110000
                ;mem[7448] <= 30'b000000010000000000010110000000
                ;mem[7449] <= 30'b000000010000000000011010010000
                ;mem[7450] <= 30'b000000010000000000011010100000
                ;mem[7451] <= 30'b000000010000000000011010110000
                ;mem[7452] <= 30'b000000010000000000011100110000
                ;mem[7453] <= 30'b000000010000000000011101000000
                ;mem[7454] <= 30'b000000010000000000100001010000
                ;mem[7455] <= 30'b000000010000000000100001100000
                ;mem[7456] <= 30'b000000010000000000100001110000
                ;mem[7457] <= 30'b000000010000000000100011110000
                ;mem[7458] <= 30'b000000010000000000100100000000
                ;mem[7459] <= 30'b000000010000000000101000010000
                ;mem[7460] <= 30'b000000010000000000101000100000
                ;mem[7461] <= 30'b000000010000000000101010100000
                ;mem[7462] <= 30'b000000010000000000101010110000
                ;mem[7463] <= 30'b000000010000000000101111010000
                ;mem[7464] <= 30'b000000010000000000101111100000
                ;mem[7465] <= 30'b000000010000000000110001100000
                ;mem[7466] <= 30'b000000010000000000110001110000
                ;mem[7467] <= 30'b000000010000000000110110010000
                ;mem[7468] <= 30'b000000010000000000110110100000
                ;mem[7469] <= 30'b000000010000000000110110110000
                ;mem[7470] <= 30'b000000010000000000111000010000
                ;mem[7471] <= 30'b000000010000000000111000100000
                ;mem[7472] <= 30'b000000010000000000111000110000
                ;mem[7473] <= 30'b000000010000000000111101010000
                ;mem[7474] <= 30'b000000010000000000111101100000
                ;mem[7475] <= 30'b000000010000000000111101110000
                ;mem[7476] <= 30'b000000010000000000111111000000
                ;mem[7477] <= 30'b000000010000000000111111010000
                ;mem[7478] <= 30'b000000010000000000111111100000
                ;mem[7479] <= 30'b000000000000000001000011010000
                ;mem[7480] <= 30'b000000000000000001000011100000
                ;mem[7481] <= 30'b000000000000000001000101100000
                ;mem[7482] <= 30'b000000000000000001000101110000
                ;mem[7483] <= 30'b000000000000000001001010010000
                ;mem[7484] <= 30'b000000000000000001001010100000
                ;mem[7485] <= 30'b000000000000000001001010110000
                ;mem[7486] <= 30'b000000000000000001001100010000
                ;mem[7487] <= 30'b000000000000000001001100100000
                ;mem[7488] <= 30'b000000000000000001001100110000
                ;mem[7489] <= 30'b000000000000000001010001010000
                ;mem[7490] <= 30'b000000000000000001010001100000
                ;mem[7491] <= 30'b000000000000000001010001110000
                ;mem[7492] <= 30'b000000000000000001010011000000
                ;mem[7493] <= 30'b000000000000000001010011010000
                ;mem[7494] <= 30'b000000000000000001010011100000
                ;mem[7495] <= 30'b000000000000000001011000100000
                ;mem[7496] <= 30'b000000000000000001011000110000
                ;mem[7497] <= 30'b000000000000000001011001000000
                ;mem[7498] <= 30'b000000000000000001011001010000
                ;mem[7499] <= 30'b000000000000000001011001100000
                ;mem[7500] <= 30'b000000000000000001011001110000
                ;mem[7501] <= 30'b000000000000000001011010000000
                ;mem[7502] <= 30'b000000000000000001011010010000
                ;mem[7503] <= 30'b000000000000000001011111100000
                ;mem[7504] <= 30'b000000000000000001011111110000
                ;mem[7505] <= 30'b000000000000000001100000000000
                ;mem[7506] <= 30'b000000000000000001100000010000
                ;mem[7507] <= 30'b000000000000000001100000100000
                ;mem[7508] <= 30'b000000000000000001100000110000
                ;mem[7509] <= 30'b000000000000000001100001000000
                ;mem[7510] <= 30'b000000000000000001100111000000
                ;mem[7511] <= 30'b000000000000000001100111010000
                ;mem[7512] <= 30'b000000000000000001100111100000
                ;mem[7513] <= 30'b000000000000000000100101010000
                ;mem[7514] <= 30'b000000000000000000100101100000
                ;mem[7515] <= 30'b000000000000000000101100000000
                ;mem[7516] <= 30'b000000000000000000101100010000
                ;mem[7517] <= 30'b000000000000000000101100100000
                ;mem[7518] <= 30'b000000000000000000101111000000
                ;mem[7519] <= 30'b000000000000000000101111010000
                ;mem[7520] <= 30'b000000000000000000110011000000
                ;mem[7521] <= 30'b000000000000000000110011010000
                ;mem[7522] <= 30'b000000000000000000110011100000
                ;mem[7523] <= 30'b000000000000000000110110000000
                ;mem[7524] <= 30'b000000000000000000110110010000
                ;mem[7525] <= 30'b000000000000000000110110100000
                ;mem[7526] <= 30'b000000000000000000111010000000
                ;mem[7527] <= 30'b000000000000000000111010010000
                ;mem[7528] <= 30'b000000000000000000111010100000
                ;mem[7529] <= 30'b000000000000000000111100110000
                ;mem[7530] <= 30'b000000000000000000111101000000
                ;mem[7531] <= 30'b000000000000000000111101010000
                ;mem[7532] <= 30'b000000001000000000000000000000
                ;mem[7533] <= 30'b000000001000000000000000010000
                ;mem[7534] <= 30'b000000001000000000000000100000
                ;mem[7535] <= 30'b000000001000000000000011000000
                ;mem[7536] <= 30'b000000001000000000000011010000
                ;mem[7537] <= 30'b000000001000000000000111000000
                ;mem[7538] <= 30'b000000001000000000000111010000
                ;mem[7539] <= 30'b000000001000000000000111100000
                ;mem[7540] <= 30'b000000001000000000001010000000
                ;mem[7541] <= 30'b000000001000000000001010010000
                ;mem[7542] <= 30'b000000001000000000001010100000
                ;mem[7543] <= 30'b000000001000000000001110000000
                ;mem[7544] <= 30'b000000001000000000001110010000
                ;mem[7545] <= 30'b000000001000000000001110100000
                ;mem[7546] <= 30'b000000001000000000010000110000
                ;mem[7547] <= 30'b000000001000000000010001000000
                ;mem[7548] <= 30'b000000001000000000010001010000
                ;mem[7549] <= 30'b000000001000000000010101000000
                ;mem[7550] <= 30'b000000001000000000010101010000
                ;mem[7551] <= 30'b000000001000000000010101100000
                ;mem[7552] <= 30'b000000001000000000010111110000
                ;mem[7553] <= 30'b000000001000000000011000000000
                ;mem[7554] <= 30'b000000001000000000011000010000
                ;mem[7555] <= 30'b000000001000000000011100000000
                ;mem[7556] <= 30'b000000001000000000011100010000
                ;mem[7557] <= 30'b000000001000000000011100100000
                ;mem[7558] <= 30'b000000001000000000011110110000
                ;mem[7559] <= 30'b000000001000000000011111000000
                ;mem[7560] <= 30'b000000001000000000011111010000
                ;mem[7561] <= 30'b000000001000000000100010110000
                ;mem[7562] <= 30'b000000001000000000100011000000
                ;mem[7563] <= 30'b000000001000000000100011010000
                ;mem[7564] <= 30'b000000001000000000100011100000
                ;mem[7565] <= 30'b000000001000000000100101110000
                ;mem[7566] <= 30'b000000001000000000100110000000
                ;mem[7567] <= 30'b000000001000000000101001110000
                ;mem[7568] <= 30'b000000001000000000101010000000
                ;mem[7569] <= 30'b000000001000000000101010010000
                ;mem[7570] <= 30'b000000001000000000101100110000
                ;mem[7571] <= 30'b000000001000000000101101000000
                ;mem[7572] <= 30'b000000001000000000110000110000
                ;mem[7573] <= 30'b000000001000000000110001000000
                ;mem[7574] <= 30'b000000001000000000110001010000
                ;mem[7575] <= 30'b000000001000000000110011100000
                ;mem[7576] <= 30'b000000001000000000110011110000
                ;mem[7577] <= 30'b000000001000000000110100000000
                ;mem[7578] <= 30'b000000001000000000110111110000
                ;mem[7579] <= 30'b000000001000000000111000000000
                ;mem[7580] <= 30'b000000001000000000111000010000
                ;mem[7581] <= 30'b000000001000000000111000100000
                ;mem[7582] <= 30'b000000001000000000111000110000
                ;mem[7583] <= 30'b000000001000000000111001000000
                ;mem[7584] <= 30'b000000001000000000111001010000
                ;mem[7585] <= 30'b000000001000000000111001100000
                ;mem[7586] <= 30'b000000001000000000111010010000
                ;mem[7587] <= 30'b000000001000000000111010100000
                ;mem[7588] <= 30'b000000001000000000111010110000
                ;mem[7589] <= 30'b000000001000000000111011000000
                ;mem[7590] <= 30'b000000001000000000111110110000
                ;mem[7591] <= 30'b000000001000000000111111000000
                ;mem[7592] <= 30'b000000001000000000111111010000
                ;mem[7593] <= 30'b000000001000000000111111100000
                ;mem[7594] <= 30'b000000001000000000111111110000
                ;mem[7595] <= 30'b000000010000000000000000110000
                ;mem[7596] <= 30'b000000010000000000000001000000
                ;mem[7597] <= 30'b000000010000000000000100110000
                ;mem[7598] <= 30'b000000010000000000000101000000
                ;mem[7599] <= 30'b000000010000000000000101010000
                ;mem[7600] <= 30'b000000010000000000000111100000
                ;mem[7601] <= 30'b000000010000000000000111110000
                ;mem[7602] <= 30'b000000010000000000001000000000
                ;mem[7603] <= 30'b000000010000000000001011110000
                ;mem[7604] <= 30'b000000010000000000001100000000
                ;mem[7605] <= 30'b000000010000000000001100010000
                ;mem[7606] <= 30'b000000010000000000001100100000
                ;mem[7607] <= 30'b000000010000000000001100110000
                ;mem[7608] <= 30'b000000010000000000001101000000
                ;mem[7609] <= 30'b000000010000000000001101010000
                ;mem[7610] <= 30'b000000010000000000001101100000
                ;mem[7611] <= 30'b000000010000000000001110010000
                ;mem[7612] <= 30'b000000010000000000001110100000
                ;mem[7613] <= 30'b000000010000000000001110110000
                ;mem[7614] <= 30'b000000010000000000001111000000
                ;mem[7615] <= 30'b000000010000000000010010110000
                ;mem[7616] <= 30'b000000010000000000010011000000
                ;mem[7617] <= 30'b000000010000000000010011010000
                ;mem[7618] <= 30'b000000010000000000010011100000
                ;mem[7619] <= 30'b000000010000000000010011110000
                ;mem[7620] <= 30'b000000010000000000010100000000
                ;mem[7621] <= 30'b000000010000000000010100010000
                ;mem[7622] <= 30'b000000010000000000010100100000
                ;mem[7623] <= 30'b000000010000000000010100110000
                ;mem[7624] <= 30'b000000010000000000010101000000
                ;mem[7625] <= 30'b000000010000000000010101010000
                ;mem[7626] <= 30'b000000010000000000010101100000
                ;mem[7627] <= 30'b000000010000000000010101110000
                ;mem[7628] <= 30'b000000010000000000010110000000
                ;mem[7629] <= 30'b000000010000000000011001110000
                ;mem[7630] <= 30'b000000010000000000011010000000
                ;mem[7631] <= 30'b000000010000000000011010010000
                ;mem[7632] <= 30'b000000010000000000011010100000
                ;mem[7633] <= 30'b000000010000000000011010110000
                ;mem[7634] <= 30'b000000010000000000011011000000
                ;mem[7635] <= 30'b000000010000000000011011010000
                ;mem[7636] <= 30'b000000010000000000011011100000
                ;mem[7637] <= 30'b000000010000000000011011110000
                ;mem[7638] <= 30'b000000010000000000011100000000
                ;mem[7639] <= 30'b000000010000000000011100010000
                ;mem[7640] <= 30'b000000010000000000011100100000
                ;mem[7641] <= 30'b000000010000000000011100110000
                ;mem[7642] <= 30'b000000010000000000011101000000
                ;mem[7643] <= 30'b000000010000000000100001000000
                ;mem[7644] <= 30'b000000010000000000100001010000
                ;mem[7645] <= 30'b000000010000000000100011010000
                ;mem[7646] <= 30'b000000010000000000100011100000
                ;mem[7647] <= 30'b000000010000000000100011110000
                ;mem[7648] <= 30'b000000010000000000101010010000
                ;mem[7649] <= 30'b000000010000000000101010100000
                ;mem[7650] <= 30'b000000010000000000110001000000
                ;mem[7651] <= 30'b000000010000000000110001010000
                ;mem[7652] <= 30'b000000010000000000110001100000
                ;mem[7653] <= 30'b000000010000000000111000000000
                ;mem[7654] <= 30'b000000010000000000111000010000
                ;mem[7655] <= 30'b000000010000000000111000100000
                ;mem[7656] <= 30'b000000010000000000111111000000
                ;mem[7657] <= 30'b000000010000000000111111010000
                ;mem[7658] <= 30'b000000010000000000111111100000
                ;mem[7659] <= 30'b000000000000000001000101000000
                ;mem[7660] <= 30'b000000000000000001000101010000
                ;mem[7661] <= 30'b000000000000000001000101100000
                ;mem[7662] <= 30'b000000000000000001001100000000
                ;mem[7663] <= 30'b000000000000000001001100010000
                ;mem[7664] <= 30'b000000000000000001001100100000
                ;mem[7665] <= 30'b000000000000000001010011000000
                ;mem[7666] <= 30'b000000000000000001010011010000
                ;mem[7667] <= 30'b000000000000000001010011100000
                ;mem[7668] <= 30'b000000000000000001011010000000
                ;mem[7669] <= 30'b000000000000000001011010010000
                ;mem[7670] <= 30'b000000000000000001011010100000
                ;mem[7671] <= 30'b000000000000000001100001000000
                ;mem[7672] <= 30'b000000000000000001100001010000
                ;mem[7673] <= 30'b000000000000000001100001100000
                ;mem[7674] <= 30'b000000000000000001101000000000
                ;mem[7675] <= 30'b000000000000000001101000010000
                ;mem[7676] <= 30'b000000000000000000100111000000
                ;mem[7677] <= 30'b000000000000000000101101110000
                ;mem[7678] <= 30'b000000000000000000101110000000
                ;mem[7679] <= 30'b000000000000000000101110010000
                ;mem[7680] <= 30'b000000000000000000110100110000
                ;mem[7681] <= 30'b000000000000000000110101000000
                ;mem[7682] <= 30'b000000000000000000110101010000
                ;mem[7683] <= 30'b000000000000000000111011110000
                ;mem[7684] <= 30'b000000000000000000111100000000
                ;mem[7685] <= 30'b000000001000000000000001110000
                ;mem[7686] <= 30'b000000001000000000000010000000
                ;mem[7687] <= 30'b000000001000000000000010010000
                ;mem[7688] <= 30'b000000001000000000001000110000
                ;mem[7689] <= 30'b000000001000000000001001000000
                ;mem[7690] <= 30'b000000001000000000001001010000
                ;mem[7691] <= 30'b000000001000000000001111110000
                ;mem[7692] <= 30'b000000001000000000010000000000
                ;mem[7693] <= 30'b000000001000000000010110110000
                ;mem[7694] <= 30'b000000001000000000010111000000
                ;mem[7695] <= 30'b000000001000000000011101110000
                ;mem[7696] <= 30'b000000001000000000011110000000
                ;mem[7697] <= 30'b000000001000000000100100100000
                ;mem[7698] <= 30'b000000001000000000100100110000
                ;mem[7699] <= 30'b000000001000000000100101000000
                ;mem[7700] <= 30'b000000001000000000101011100000
                ;mem[7701] <= 30'b000000001000000000101011110000
                ;mem[7702] <= 30'b000000001000000000110010100000
                ;mem[7703] <= 30'b000000001000000000110010110000
                ;mem[7704] <= 30'b000000001000000000111001100000
                ;mem[7705] <= 30'b000000010000000000000110100000
                ;mem[7706] <= 30'b000000010000000000000110110000
                ;mem[7707] <= 30'b000000010000000000001101100000
                ;mem[7708] <= 30'b000000010000000000010100100000
                ;mem[7709] <= 30'b000000010000000000011011010000
                ;mem[7710] <= 30'b000000010000000000011011100000
                ;mem[7711] <= 30'b000000010000000000100010010000
                ;mem[7712] <= 30'b000000010000000000100010100000
                ;mem[7713] <= 30'b000000010000000000101001000000
                ;mem[7714] <= 30'b000000010000000000101001010000
                ;mem[7715] <= 30'b000000010000000000110000000000
                ;mem[7716] <= 30'b000000010000000000110000010000
                ;mem[7717] <= 30'b000000010000000000110111000000
                ;mem[7718] <= 30'b000000010000000000110111010000
                ;mem[7719] <= 30'b000000010000000000111110000000
                ;mem[7720] <= 30'b000000010000000000111110010000
                ;mem[7721] <= 30'b000000000000000001000100000000
                ;mem[7722] <= 30'b000000000000000001000100010000
                ;mem[7723] <= 30'b000000000000000001001011000000
                ;mem[7724] <= 30'b000000000000000001001011010000
                ;mem[7725] <= 30'b000000000000000001010010000000
                ;mem[7726] <= 30'b000000000000000001010010010000
                ;mem[7727] <= 30'b000000000000000001011001000000
                ;mem[7728] <= 30'b000000000000000001011001010000
                ;mem[7729] <= 30'b000000000000000001100000000000
                ;mem[7730] <= 30'b000000000000000001100000010000
                ;mem[7731] <= 30'b000000000000000001100111000000
                ;mem[7732] <= 30'b000000000000000001100111010000
                ;mem[7733] <= 30'b000000000000000000110100110000
                ;mem[7734] <= 30'b000000000000000000110101000000
                ;mem[7735] <= 30'b000000000000000000110101010000
                ;mem[7736] <= 30'b000000000000000000110101100000
                ;mem[7737] <= 30'b000000000000000000111011000000
                ;mem[7738] <= 30'b000000000000000000111011010000
                ;mem[7739] <= 30'b000000000000000000111011100000
                ;mem[7740] <= 30'b000000000000000000111011110000
                ;mem[7741] <= 30'b000000000000000000111100000000
                ;mem[7742] <= 30'b000000000000000000111100010000
                ;mem[7743] <= 30'b000000000000000000111100100000
                ;mem[7744] <= 30'b000000000000000000111100110000
                ;mem[7745] <= 30'b000000001000000000001000110000
                ;mem[7746] <= 30'b000000001000000000001001000000
                ;mem[7747] <= 30'b000000001000000000001001010000
                ;mem[7748] <= 30'b000000001000000000001001100000
                ;mem[7749] <= 30'b000000001000000000001111000000
                ;mem[7750] <= 30'b000000001000000000001111010000
                ;mem[7751] <= 30'b000000001000000000001111100000
                ;mem[7752] <= 30'b000000001000000000001111110000
                ;mem[7753] <= 30'b000000001000000000010000000000
                ;mem[7754] <= 30'b000000001000000000010000010000
                ;mem[7755] <= 30'b000000001000000000010000100000
                ;mem[7756] <= 30'b000000001000000000010000110000
                ;mem[7757] <= 30'b000000001000000000010101100000
                ;mem[7758] <= 30'b000000001000000000010101110000
                ;mem[7759] <= 30'b000000001000000000010110000000
                ;mem[7760] <= 30'b000000001000000000010110010000
                ;mem[7761] <= 30'b000000001000000000010110100000
                ;mem[7762] <= 30'b000000001000000000010110110000
                ;mem[7763] <= 30'b000000001000000000010111010000
                ;mem[7764] <= 30'b000000001000000000010111100000
                ;mem[7765] <= 30'b000000001000000000010111110000
                ;mem[7766] <= 30'b000000001000000000011100010000
                ;mem[7767] <= 30'b000000001000000000011100100000
                ;mem[7768] <= 30'b000000001000000000011100110000
                ;mem[7769] <= 30'b000000001000000000011101000000
                ;mem[7770] <= 30'b000000001000000000011110100000
                ;mem[7771] <= 30'b000000001000000000011110110000
                ;mem[7772] <= 30'b000000001000000000100011000000
                ;mem[7773] <= 30'b000000001000000000100011010000
                ;mem[7774] <= 30'b000000001000000000100011100000
                ;mem[7775] <= 30'b000000001000000000100101100000
                ;mem[7776] <= 30'b000000001000000000100101110000
                ;mem[7777] <= 30'b000000001000000000100110000000
                ;mem[7778] <= 30'b000000001000000000101001110000
                ;mem[7779] <= 30'b000000001000000000101010000000
                ;mem[7780] <= 30'b000000001000000000101010010000
                ;mem[7781] <= 30'b000000001000000000101100100000
                ;mem[7782] <= 30'b000000001000000000101100110000
                ;mem[7783] <= 30'b000000001000000000101101000000
                ;mem[7784] <= 30'b000000001000000000110000100000
                ;mem[7785] <= 30'b000000001000000000110000110000
                ;mem[7786] <= 30'b000000001000000000110001000000
                ;mem[7787] <= 30'b000000001000000000110011010000
                ;mem[7788] <= 30'b000000001000000000110011100000
                ;mem[7789] <= 30'b000000001000000000110011110000
                ;mem[7790] <= 30'b000000001000000000110100000000
                ;mem[7791] <= 30'b000000001000000000110111100000
                ;mem[7792] <= 30'b000000001000000000110111110000
                ;mem[7793] <= 30'b000000001000000000111000000000
                ;mem[7794] <= 30'b000000001000000000111001100000
                ;mem[7795] <= 30'b000000001000000000111001110000
                ;mem[7796] <= 30'b000000001000000000111010000000
                ;mem[7797] <= 30'b000000001000000000111010010000
                ;mem[7798] <= 30'b000000001000000000111010100000
                ;mem[7799] <= 30'b000000001000000000111010110000
                ;mem[7800] <= 30'b000000001000000000111011000000
                ;mem[7801] <= 30'b000000001000000000111110110000
                ;mem[7802] <= 30'b000000001000000000111111000000
                ;mem[7803] <= 30'b000000001000000000111111010000
                ;mem[7804] <= 30'b000000001000000000111111100000
                ;mem[7805] <= 30'b000000001000000000111111110000
                ;mem[7806] <= 30'b000000010000000000000000100000
                ;mem[7807] <= 30'b000000010000000000000000110000
                ;mem[7808] <= 30'b000000010000000000000001000000
                ;mem[7809] <= 30'b000000010000000000000100100000
                ;mem[7810] <= 30'b000000010000000000000100110000
                ;mem[7811] <= 30'b000000010000000000000101000000
                ;mem[7812] <= 30'b000000010000000000000111010000
                ;mem[7813] <= 30'b000000010000000000000111100000
                ;mem[7814] <= 30'b000000010000000000000111110000
                ;mem[7815] <= 30'b000000010000000000001000000000
                ;mem[7816] <= 30'b000000010000000000001011100000
                ;mem[7817] <= 30'b000000010000000000001011110000
                ;mem[7818] <= 30'b000000010000000000001100000000
                ;mem[7819] <= 30'b000000010000000000001101100000
                ;mem[7820] <= 30'b000000010000000000001101110000
                ;mem[7821] <= 30'b000000010000000000001110000000
                ;mem[7822] <= 30'b000000010000000000001110010000
                ;mem[7823] <= 30'b000000010000000000001110100000
                ;mem[7824] <= 30'b000000010000000000001110110000
                ;mem[7825] <= 30'b000000010000000000001111000000
                ;mem[7826] <= 30'b000000010000000000010010110000
                ;mem[7827] <= 30'b000000010000000000010011000000
                ;mem[7828] <= 30'b000000010000000000010011010000
                ;mem[7829] <= 30'b000000010000000000010011100000
                ;mem[7830] <= 30'b000000010000000000010011110000
                ;mem[7831] <= 30'b000000010000000000010100000000
                ;mem[7832] <= 30'b000000010000000000010100010000
                ;mem[7833] <= 30'b000000010000000000010100100000
                ;mem[7834] <= 30'b000000010000000000010100110000
                ;mem[7835] <= 30'b000000010000000000010101000000
                ;mem[7836] <= 30'b000000010000000000010101010000
                ;mem[7837] <= 30'b000000010000000000010101100000
                ;mem[7838] <= 30'b000000010000000000010101110000
                ;mem[7839] <= 30'b000000010000000000011010000000
                ;mem[7840] <= 30'b000000010000000000011010010000
                ;mem[7841] <= 30'b000000010000000000011010100000
                ;mem[7842] <= 30'b000000010000000000011010110000
                ;mem[7843] <= 30'b000000010000000000011011000000
                ;mem[7844] <= 30'b000000010000000000011011010000
                ;mem[7845] <= 30'b000000010000000000011011100000
                ;mem[7846] <= 30'b000000010000000000011100010000
                ;mem[7847] <= 30'b000000010000000000011100100000
                ;mem[7848] <= 30'b000000010000000000011100110000
                ;mem[7849] <= 30'b000000010000000000100011010000
                ;mem[7850] <= 30'b000000010000000000100011100000
                ;mem[7851] <= 30'b000000010000000000101010000000
                ;mem[7852] <= 30'b000000010000000000101010010000
                ;mem[7853] <= 30'b000000010000000000101010100000
                ;mem[7854] <= 30'b000000010000000000110001000000
                ;mem[7855] <= 30'b000000010000000000110001010000
                ;mem[7856] <= 30'b000000010000000000111000000000
                ;mem[7857] <= 30'b000000010000000000111000010000
                ;mem[7858] <= 30'b000000010000000000111110110000
                ;mem[7859] <= 30'b000000010000000000111111000000
                ;mem[7860] <= 30'b000000010000000000111111010000
                ;mem[7861] <= 30'b000000000000000001000101000000
                ;mem[7862] <= 30'b000000000000000001000101010000
                ;mem[7863] <= 30'b000000000000000001001100000000
                ;mem[7864] <= 30'b000000000000000001001100010000
                ;mem[7865] <= 30'b000000000000000001010010110000
                ;mem[7866] <= 30'b000000000000000001010011000000
                ;mem[7867] <= 30'b000000000000000001010011010000
                ;mem[7868] <= 30'b000000000000000001011001110000
                ;mem[7869] <= 30'b000000000000000001011010000000
                ;mem[7870] <= 30'b000000000000000001011010010000
                ;mem[7871] <= 30'b000000000000000001100000100000
                ;mem[7872] <= 30'b000000000000000001100000110000
                ;mem[7873] <= 30'b000000000000000001100001000000
                ;mem[7874] <= 30'b000000000000000001100111100000
                ;mem[7875] <= 30'b000000000000000001100111110000
                ;mem[7876] <= 30'b000000000000000001101000000000
                ;mem[7877] <= 30'b000000000000000001101110010000
                ;mem[7878] <= 30'b000000000000000001101110100000
                ;mem[7879] <= 30'b000000000000000001101110110000
                ;mem[7880] <= 30'b000000000000000001110101100000
                ;mem[7881] <= 30'b000000000000000000110000000000
                ;mem[7882] <= 30'b000000000000000000110110100000
                ;mem[7883] <= 30'b000000000000000000110110110000
                ;mem[7884] <= 30'b000000000000000000111100100000
                ;mem[7885] <= 30'b000000000000000000111100110000
                ;mem[7886] <= 30'b000000000000000000111101000000
                ;mem[7887] <= 30'b000000000000000000111101010000
                ;mem[7888] <= 30'b000000001000000000000100000000
                ;mem[7889] <= 30'b000000001000000000001010100000
                ;mem[7890] <= 30'b000000001000000000001010110000
                ;mem[7891] <= 30'b000000001000000000010000100000
                ;mem[7892] <= 30'b000000001000000000010000110000
                ;mem[7893] <= 30'b000000001000000000010001000000
                ;mem[7894] <= 30'b000000001000000000010001010000
                ;mem[7895] <= 30'b000000001000000000010110110000
                ;mem[7896] <= 30'b000000001000000000010111000000
                ;mem[7897] <= 30'b000000001000000000010111010000
                ;mem[7898] <= 30'b000000001000000000010111100000
                ;mem[7899] <= 30'b000000001000000000010111110000
                ;mem[7900] <= 30'b000000001000000000011100110000
                ;mem[7901] <= 30'b000000001000000000011101000000
                ;mem[7902] <= 30'b000000001000000000011101010000
                ;mem[7903] <= 30'b000000001000000000011101100000
                ;mem[7904] <= 30'b000000001000000000011101110000
                ;mem[7905] <= 30'b000000001000000000011110000000
                ;mem[7906] <= 30'b000000001000000000011110010000
                ;mem[7907] <= 30'b000000001000000000100011100000
                ;mem[7908] <= 30'b000000001000000000100011110000
                ;mem[7909] <= 30'b000000001000000000100100000000
                ;mem[7910] <= 30'b000000001000000000100100010000
                ;mem[7911] <= 30'b000000001000000000100100100000
                ;mem[7912] <= 30'b000000001000000000111000010000
                ;mem[7913] <= 30'b000000001000000000111111010000
                ;mem[7914] <= 30'b000000001000000000111111100000
                ;mem[7915] <= 30'b000000010000000000001100010000
                ;mem[7916] <= 30'b000000010000000000010011010000
                ;mem[7917] <= 30'b000000010000000000010011100000
                ;mem[7918] <= 30'b000000010000000000011010010000
                ;mem[7919] <= 30'b000000010000000000011010100000
                ;mem[7920] <= 30'b000000010000000000011010110000
                ;mem[7921] <= 30'b000000010000000000011011000000
                ;mem[7922] <= 30'b000000010000000000100010000000
                ;mem[7923] <= 30'b000000010000000000100010010000
                ;mem[7924] <= 30'b000000010000000000101001000000
                ;mem[7925] <= 30'b000000010000000000101001010000
                ;mem[7926] <= 30'b000000010000000000110000000000
                ;mem[7927] <= 30'b000000010000000000110000010000
                ;mem[7928] <= 30'b000000010000000000110111000000
                ;mem[7929] <= 30'b000000010000000000111110000000
                ;mem[7930] <= 30'b000000000000000001000100000000
                ;mem[7931] <= 30'b000000000000000001000100010000
                ;mem[7932] <= 30'b000000000000000001001011000000
                ;mem[7933] <= 30'b000000000000000001010010000000
                ;mem[7934] <= 30'b000000000000000001011000110000
                ;mem[7935] <= 30'b000000000000000001011001000000
                ;mem[7936] <= 30'b000000000000000001011111110000
                ;mem[7937] <= 30'b000000000000000001100000000000
                ;mem[7938] <= 30'b000000000000000001100110100000
                ;mem[7939] <= 30'b000000000000000001100110110000
                ;mem[7940] <= 30'b000000000000000001101101100000
                ;mem[7941] <= 30'b000000000000000000110001110000
                ;mem[7942] <= 30'b000000000000000000110010000000
                ;mem[7943] <= 30'b000000000000000000110010010000
                ;mem[7944] <= 30'b000000000000000000110010100000
                ;mem[7945] <= 30'b000000000000000000110010110000
                ;mem[7946] <= 30'b000000000000000000111000100000
                ;mem[7947] <= 30'b000000000000000000111000110000
                ;mem[7948] <= 30'b000000000000000000111001000000
                ;mem[7949] <= 30'b000000000000000000111001010000
                ;mem[7950] <= 30'b000000000000000000111001100000
                ;mem[7951] <= 30'b000000000000000000111001110000
                ;mem[7952] <= 30'b000000000000000000111010000000
                ;mem[7953] <= 30'b000000000000000000111010010000
                ;mem[7954] <= 30'b000000000000000000111010100000
                ;mem[7955] <= 30'b000000000000000000111010110000
                ;mem[7956] <= 30'b000000000000000000111011000000
                ;mem[7957] <= 30'b000000000000000000111011010000
                ;mem[7958] <= 30'b000000000000000000111011100000
                ;mem[7959] <= 30'b000000000000000000111111110000
                ;mem[7960] <= 30'b000000001000000000000101110000
                ;mem[7961] <= 30'b000000001000000000000110000000
                ;mem[7962] <= 30'b000000001000000000000110010000
                ;mem[7963] <= 30'b000000001000000000000110100000
                ;mem[7964] <= 30'b000000001000000000000110110000
                ;mem[7965] <= 30'b000000001000000000001100100000
                ;mem[7966] <= 30'b000000001000000000001100110000
                ;mem[7967] <= 30'b000000001000000000001101000000
                ;mem[7968] <= 30'b000000001000000000001101010000
                ;mem[7969] <= 30'b000000001000000000001101100000
                ;mem[7970] <= 30'b000000001000000000001101110000
                ;mem[7971] <= 30'b000000001000000000001110000000
                ;mem[7972] <= 30'b000000001000000000001110010000
                ;mem[7973] <= 30'b000000001000000000001110100000
                ;mem[7974] <= 30'b000000001000000000001110110000
                ;mem[7975] <= 30'b000000001000000000001111000000
                ;mem[7976] <= 30'b000000001000000000001111010000
                ;mem[7977] <= 30'b000000001000000000001111100000
                ;mem[7978] <= 30'b000000001000000000010011110000
                ;mem[7979] <= 30'b000000001000000000010100000000
                ;mem[7980] <= 30'b000000001000000000010100010000
                ;mem[7981] <= 30'b000000001000000000010100100000
                ;mem[7982] <= 30'b000000001000000000010100110000
                ;mem[7983] <= 30'b000000001000000000010101000000
                ;mem[7984] <= 30'b000000001000000000010101010000
                ;mem[7985] <= 30'b000000001000000000010101100000
                ;mem[7986] <= 30'b000000001000000000010101110000
                ;mem[7987] <= 30'b000000001000000000010110000000
                ;mem[7988] <= 30'b000000001000000000010110010000
                ;mem[7989] <= 30'b000000001000000000010110100000
                ;mem[7990] <= 30'b000000001000000000010110110000
                ;mem[7991] <= 30'b000000001000000000010111000000
                ;mem[7992] <= 30'b000000001000000000011011100000
                ;mem[7993] <= 30'b000000001000000000011011110000
                ;mem[7994] <= 30'b000000001000000000011100000000
                ;mem[7995] <= 30'b000000001000000000011100010000
                ;mem[7996] <= 30'b000000001000000000011100100000
                ;mem[7997] <= 30'b000000001000000000011100110000
                ;mem[7998] <= 30'b000000001000000000011101000000
                ;mem[7999] <= 30'b000000001000000000011101010000
                ;mem[8000] <= 30'b000000001000000000011101100000
                ;mem[8001] <= 30'b000000001000000000011101110000
                ;mem[8002] <= 30'b000000001000000000011110000000
                ;mem[8003] <= 30'b000000001000000000011110010000
                ;mem[8004] <= 30'b000000001000000000011110100000
                ;mem[8005] <= 30'b000000001000000000100100100000
                ;mem[8006] <= 30'b000000001000000000100100110000
                ;mem[8007] <= 30'b000000001000000000100101000000
                ;mem[8008] <= 30'b000000001000000000100101010000
                ;mem[8009] <= 30'b000000001000000000100101100000
                ;mem[8010] <= 30'b000000001000000000100101110000
                ;mem[8011] <= 30'b000000001000000000101100000000
                ;mem[8012] <= 30'b000000001000000000101100010000
                ;mem[8013] <= 30'b000000001000000000101100100000
                ;mem[8014] <= 30'b000000001000000000101100110000
                ;mem[8015] <= 30'b000000001000000000101101000000
                ;mem[8016] <= 30'b000000001000000000110011010000
                ;mem[8017] <= 30'b000000001000000000110011100000
                ;mem[8018] <= 30'b000000001000000000110011110000
                ;mem[8019] <= 30'b000000001000000000110100000000
                ;mem[8020] <= 30'b000000001000000000111010010000
                ;mem[8021] <= 30'b000000001000000000111010100000
                ;mem[8022] <= 30'b000000001000000000111010110000
                ;mem[8023] <= 30'b000000001000000000111011000000
                ;mem[8024] <= 30'b000000010000000000000000000000
                ;mem[8025] <= 30'b000000010000000000000000010000
                ;mem[8026] <= 30'b000000010000000000000000100000
                ;mem[8027] <= 30'b000000010000000000000000110000
                ;mem[8028] <= 30'b000000010000000000000001000000
                ;mem[8029] <= 30'b000000010000000000000111010000
                ;mem[8030] <= 30'b000000010000000000000111100000
                ;mem[8031] <= 30'b000000010000000000000111110000
                ;mem[8032] <= 30'b000000010000000000001000000000
                ;mem[8033] <= 30'b000000010000000000001110010000
                ;mem[8034] <= 30'b000000010000000000001110100000
                ;mem[8035] <= 30'b000000010000000000001110110000
                ;mem[8036] <= 30'b000000010000000000001111000000
                ;mem[8037] <= 30'b000000010000000000010101010000
                ;mem[8038] <= 30'b000000010000000000010101100000
                ;mem[8039] <= 30'b000000010000000000010101110000
                ;mem[8040] <= 30'b000000010000000000010110000000
                ;mem[8041] <= 30'b000000010000000000011100010000
                ;mem[8042] <= 30'b000000010000000000011100100000
                ;mem[8043] <= 30'b000000010000000000011100110000
                ;mem[8044] <= 30'b000000010000000000011101000000
                ;mem[8045] <= 30'b000000010000000000011101010000
                ;mem[8046] <= 30'b000000010000000000100011010000
                ;mem[8047] <= 30'b000000010000000000100011100000
                ;mem[8048] <= 30'b000000010000000000100011110000
                ;mem[8049] <= 30'b000000010000000000100100000000
                ;mem[8050] <= 30'b000000010000000000101010010000
                ;mem[8051] <= 30'b000000010000000000101010100000
                ;mem[8052] <= 30'b000000010000000000101010110000
                ;mem[8053] <= 30'b000000010000000000101011000000
                ;mem[8054] <= 30'b000000010000000000110001010000
                ;mem[8055] <= 30'b000000010000000000110001100000
                ;mem[8056] <= 30'b000000010000000000110001110000
                ;mem[8057] <= 30'b000000010000000000110010000000
                ;mem[8058] <= 30'b000000010000000000111000000000
                ;mem[8059] <= 30'b000000010000000000111000010000
                ;mem[8060] <= 30'b000000010000000000111000100000
                ;mem[8061] <= 30'b000000010000000000111000110000
                ;mem[8062] <= 30'b000000010000000000111111000000
                ;mem[8063] <= 30'b000000010000000000111111010000
                ;mem[8064] <= 30'b000000010000000000111111100000
                ;mem[8065] <= 30'b000000010000000000111111110000
                ;mem[8066] <= 30'b000000000000000001000101010000
                ;mem[8067] <= 30'b000000000000000001000101100000
                ;mem[8068] <= 30'b000000000000000001000101110000
                ;mem[8069] <= 30'b000000000000000001000110000000
                ;mem[8070] <= 30'b000000000000000001001100000000
                ;mem[8071] <= 30'b000000000000000001001100010000
                ;mem[8072] <= 30'b000000000000000001001100100000
                ;mem[8073] <= 30'b000000000000000001001100110000
                ;mem[8074] <= 30'b000000000000000001010011000000
                ;mem[8075] <= 30'b000000000000000001010011010000
                ;mem[8076] <= 30'b000000000000000001010011100000
                ;mem[8077] <= 30'b000000000000000001010011110000
                ;mem[8078] <= 30'b000000000000000001011010000000
                ;mem[8079] <= 30'b000000000000000001011010010000
                ;mem[8080] <= 30'b000000000000000001011010100000
                ;mem[8081] <= 30'b000000000000000001100000110000
                ;mem[8082] <= 30'b000000000000000001100001000000
                ;mem[8083] <= 30'b000000000000000001100001010000
                ;mem[8084] <= 30'b000000000000000001100001100000
                ;mem[8085] <= 30'b000000000000000001100111100000
                ;mem[8086] <= 30'b000000000000000001100111110000
                ;mem[8087] <= 30'b000000000000000001101000000000
                ;mem[8088] <= 30'b000000000000000001101000010000
                ;mem[8089] <= 30'b000000000000000001101000100000
                ;mem[8090] <= 30'b000000000000000001101110100000
                ;mem[8091] <= 30'b000000000000000001101110110000
                ;mem[8092] <= 30'b000000000000000001101111000000
                ;mem[8093] <= 30'b000000000000000001101111010000
                ;mem[8094] <= 30'b000000000000000001110101100000
                ;mem[8095] <= 30'b000000000000000001110101110000
                ;mem[8096] <= 30'b000000000000000001110110000000
                ;mem[8097] <= 30'b000000000000000000101101010000
                ;mem[8098] <= 30'b000000000000000000101101100000
                ;mem[8099] <= 30'b000000000000000000101101110000
                ;mem[8100] <= 30'b000000000000000000101110000000
                ;mem[8101] <= 30'b000000000000000000101110010000
                ;mem[8102] <= 30'b000000000000000000101110100000
                ;mem[8103] <= 30'b000000000000000000101110110000
                ;mem[8104] <= 30'b000000000000000000101111000000
                ;mem[8105] <= 30'b000000000000000000110011110000
                ;mem[8106] <= 30'b000000000000000000110100000000
                ;mem[8107] <= 30'b000000000000000000110100010000
                ;mem[8108] <= 30'b000000000000000000110100100000
                ;mem[8109] <= 30'b000000000000000000110100110000
                ;mem[8110] <= 30'b000000000000000000110101000000
                ;mem[8111] <= 30'b000000000000000000110101010000
                ;mem[8112] <= 30'b000000000000000000110101100000
                ;mem[8113] <= 30'b000000000000000000110101110000
                ;mem[8114] <= 30'b000000000000000000110110000000
                ;mem[8115] <= 30'b000000000000000000110110010000
                ;mem[8116] <= 30'b000000000000000000110110100000
                ;mem[8117] <= 30'b000000000000000000111010100000
                ;mem[8118] <= 30'b000000000000000000111010110000
                ;mem[8119] <= 30'b000000000000000000111011000000
                ;mem[8120] <= 30'b000000000000000000111011010000
                ;mem[8121] <= 30'b000000000000000000111101000000
                ;mem[8122] <= 30'b000000000000000000111101010000
                ;mem[8123] <= 30'b000000000000000000111101100000
                ;mem[8124] <= 30'b000000000000000000111101110000
                ;mem[8125] <= 30'b000000001000000000000001010000
                ;mem[8126] <= 30'b000000001000000000000001100000
                ;mem[8127] <= 30'b000000001000000000000001110000
                ;mem[8128] <= 30'b000000001000000000000010000000
                ;mem[8129] <= 30'b000000001000000000000010010000
                ;mem[8130] <= 30'b000000001000000000000010100000
                ;mem[8131] <= 30'b000000001000000000000010110000
                ;mem[8132] <= 30'b000000001000000000000011000000
                ;mem[8133] <= 30'b000000001000000000000111110000
                ;mem[8134] <= 30'b000000001000000000001000000000
                ;mem[8135] <= 30'b000000001000000000001000010000
                ;mem[8136] <= 30'b000000001000000000001000100000
                ;mem[8137] <= 30'b000000001000000000001000110000
                ;mem[8138] <= 30'b000000001000000000001001000000
                ;mem[8139] <= 30'b000000001000000000001001010000
                ;mem[8140] <= 30'b000000001000000000001001100000
                ;mem[8141] <= 30'b000000001000000000001001110000
                ;mem[8142] <= 30'b000000001000000000001010000000
                ;mem[8143] <= 30'b000000001000000000001010010000
                ;mem[8144] <= 30'b000000001000000000001010100000
                ;mem[8145] <= 30'b000000001000000000001110100000
                ;mem[8146] <= 30'b000000001000000000001110110000
                ;mem[8147] <= 30'b000000001000000000001111000000
                ;mem[8148] <= 30'b000000001000000000001111010000
                ;mem[8149] <= 30'b000000001000000000010001000000
                ;mem[8150] <= 30'b000000001000000000010001010000
                ;mem[8151] <= 30'b000000001000000000010001100000
                ;mem[8152] <= 30'b000000001000000000010001110000
                ;mem[8153] <= 30'b000000001000000000010101010000
                ;mem[8154] <= 30'b000000001000000000010101100000
                ;mem[8155] <= 30'b000000001000000000010101110000
                ;mem[8156] <= 30'b000000001000000000010110000000
                ;mem[8157] <= 30'b000000001000000000011000010000
                ;mem[8158] <= 30'b000000001000000000011000100000
                ;mem[8159] <= 30'b000000001000000000011000110000
                ;mem[8160] <= 30'b000000001000000000011100010000
                ;mem[8161] <= 30'b000000001000000000011100100000
                ;mem[8162] <= 30'b000000001000000000011100110000
                ;mem[8163] <= 30'b000000001000000000011111010000
                ;mem[8164] <= 30'b000000001000000000011111100000
                ;mem[8165] <= 30'b000000001000000000011111110000
                ;mem[8166] <= 30'b000000001000000000100011100000
                ;mem[8167] <= 30'b000000001000000000100011110000
                ;mem[8168] <= 30'b000000001000000000100110000000
                ;mem[8169] <= 30'b000000001000000000100110010000
                ;mem[8170] <= 30'b000000001000000000100110100000
                ;mem[8171] <= 30'b000000001000000000100110110000
                ;mem[8172] <= 30'b000000001000000000101010100000
                ;mem[8173] <= 30'b000000001000000000101010110000
                ;mem[8174] <= 30'b000000001000000000101011000000
                ;mem[8175] <= 30'b000000001000000000101100100000
                ;mem[8176] <= 30'b000000001000000000101100110000
                ;mem[8177] <= 30'b000000001000000000101101000000
                ;mem[8178] <= 30'b000000001000000000101101010000
                ;mem[8179] <= 30'b000000001000000000101101100000
                ;mem[8180] <= 30'b000000001000000000110001110000
                ;mem[8181] <= 30'b000000001000000000110010000000
                ;mem[8182] <= 30'b000000001000000000110010010000
                ;mem[8183] <= 30'b000000001000000000110011010000
                ;mem[8184] <= 30'b000000001000000000110011100000
                ;mem[8185] <= 30'b000000001000000000110011110000
                ;mem[8186] <= 30'b000000001000000000110100000000
                ;mem[8187] <= 30'b000000001000000000110100010000
                ;mem[8188] <= 30'b000000001000000000111001000000
                ;mem[8189] <= 30'b000000001000000000111001010000
                ;mem[8190] <= 30'b000000001000000000111001100000
                ;mem[8191] <= 30'b000000001000000000111001110000
                ;mem[8192] <= 30'b000000001000000000111010000000
                ;mem[8193] <= 30'b000000001000000000111010010000
                ;mem[8194] <= 30'b000000001000000000111010100000
                ;mem[8195] <= 30'b000000001000000000111010110000
                ;mem[8196] <= 30'b000000010000000000000000100000
                ;mem[8197] <= 30'b000000010000000000000000110000
                ;mem[8198] <= 30'b000000010000000000000001000000
                ;mem[8199] <= 30'b000000010000000000000001010000
                ;mem[8200] <= 30'b000000010000000000000001100000
                ;mem[8201] <= 30'b000000010000000000000101110000
                ;mem[8202] <= 30'b000000010000000000000110000000
                ;mem[8203] <= 30'b000000010000000000000110010000
                ;mem[8204] <= 30'b000000010000000000000111010000
                ;mem[8205] <= 30'b000000010000000000000111100000
                ;mem[8206] <= 30'b000000010000000000000111110000
                ;mem[8207] <= 30'b000000010000000000001000000000
                ;mem[8208] <= 30'b000000010000000000001000010000
                ;mem[8209] <= 30'b000000010000000000001101000000
                ;mem[8210] <= 30'b000000010000000000001101010000
                ;mem[8211] <= 30'b000000010000000000001101100000
                ;mem[8212] <= 30'b000000010000000000001101110000
                ;mem[8213] <= 30'b000000010000000000001110000000
                ;mem[8214] <= 30'b000000010000000000001110010000
                ;mem[8215] <= 30'b000000010000000000001110100000
                ;mem[8216] <= 30'b000000010000000000001110110000
                ;mem[8217] <= 30'b000000010000000000010100000000
                ;mem[8218] <= 30'b000000010000000000010100010000
                ;mem[8219] <= 30'b000000010000000000010100100000
                ;mem[8220] <= 30'b000000010000000000010100110000
                ;mem[8221] <= 30'b000000010000000000010101000000
                ;mem[8222] <= 30'b000000010000000000011010010000
                ;mem[8223] <= 30'b000000010000000000011010100000
                ;mem[8224] <= 30'b000000010000000000011010110000
                ;mem[8225] <= 30'b000000010000000000011011000000
                ;mem[8226] <= 30'b000000010000000000011011010000
                ;mem[8227] <= 30'b000000010000000000011011100000
                ;mem[8228] <= 30'b000000010000000000011011110000
                ;mem[8229] <= 30'b000000010000000000100000100000
                ;mem[8230] <= 30'b000000010000000000100000110000
                ;mem[8231] <= 30'b000000010000000000100001000000
                ;mem[8232] <= 30'b000000010000000000100001010000
                ;mem[8233] <= 30'b000000010000000000100001100000
                ;mem[8234] <= 30'b000000010000000000100001110000
                ;mem[8235] <= 30'b000000010000000000100010100000
                ;mem[8236] <= 30'b000000010000000000100010110000
                ;mem[8237] <= 30'b000000010000000000100011000000
                ;mem[8238] <= 30'b000000010000000000100111000000
                ;mem[8239] <= 30'b000000010000000000100111010000
                ;mem[8240] <= 30'b000000010000000000100111100000
                ;mem[8241] <= 30'b000000010000000000100111110000
                ;mem[8242] <= 30'b000000010000000000101000000000
                ;mem[8243] <= 30'b000000010000000000101000010000
                ;mem[8244] <= 30'b000000010000000000101001100000
                ;mem[8245] <= 30'b000000010000000000101001110000
                ;mem[8246] <= 30'b000000010000000000101010000000
                ;mem[8247] <= 30'b000000010000000000101110000000
                ;mem[8248] <= 30'b000000010000000000101110010000
                ;mem[8249] <= 30'b000000010000000000101110100000
                ;mem[8250] <= 30'b000000010000000000101110110000
                ;mem[8251] <= 30'b000000010000000000101111000000
                ;mem[8252] <= 30'b000000010000000000101111110000
                ;mem[8253] <= 30'b000000010000000000110000000000
                ;mem[8254] <= 30'b000000010000000000110000010000
                ;mem[8255] <= 30'b000000010000000000110000100000
                ;mem[8256] <= 30'b000000010000000000110000110000
                ;mem[8257] <= 30'b000000010000000000110001000000
                ;mem[8258] <= 30'b000000010000000000110101010000
                ;mem[8259] <= 30'b000000010000000000110101100000
                ;mem[8260] <= 30'b000000010000000000110101110000
                ;mem[8261] <= 30'b000000010000000000110110000000
                ;mem[8262] <= 30'b000000010000000000110110010000
                ;mem[8263] <= 30'b000000010000000000110110100000
                ;mem[8264] <= 30'b000000010000000000110110110000
                ;mem[8265] <= 30'b000000010000000000110111000000
                ;mem[8266] <= 30'b000000010000000000110111010000
                ;mem[8267] <= 30'b000000010000000000110111100000
                ;mem[8268] <= 30'b000000010000000000110111110000
                ;mem[8269] <= 30'b000000010000000000111101000000
                ;mem[8270] <= 30'b000000010000000000111101010000
                ;mem[8271] <= 30'b000000010000000000111101100000
                ;mem[8272] <= 30'b000000010000000000111101110000
                ;mem[8273] <= 30'b000000010000000000111110000000
                ;mem[8274] <= 30'b000000010000000000111110010000
                ;mem[8275] <= 30'b000000000000000001000010000000
                ;mem[8276] <= 30'b000000000000000001000010010000
                ;mem[8277] <= 30'b000000000000000001000010100000
                ;mem[8278] <= 30'b000000000000000001000010110000
                ;mem[8279] <= 30'b000000000000000001000011000000
                ;mem[8280] <= 30'b000000000000000001000011110000
                ;mem[8281] <= 30'b000000000000000001000100000000
                ;mem[8282] <= 30'b000000000000000001000100010000
                ;mem[8283] <= 30'b000000000000000001000100100000
                ;mem[8284] <= 30'b000000000000000001000100110000
                ;mem[8285] <= 30'b000000000000000001000101000000
                ;mem[8286] <= 30'b000000000000000001001001010000
                ;mem[8287] <= 30'b000000000000000001001001100000
                ;mem[8288] <= 30'b000000000000000001001001110000
                ;mem[8289] <= 30'b000000000000000001001010000000
                ;mem[8290] <= 30'b000000000000000001001010010000
                ;mem[8291] <= 30'b000000000000000001001010100000
                ;mem[8292] <= 30'b000000000000000001001010110000
                ;mem[8293] <= 30'b000000000000000001001011000000
                ;mem[8294] <= 30'b000000000000000001001011010000
                ;mem[8295] <= 30'b000000000000000001001011100000
                ;mem[8296] <= 30'b000000000000000001001011110000
                ;mem[8297] <= 30'b000000000000000001010001000000
                ;mem[8298] <= 30'b000000000000000001010001010000
                ;mem[8299] <= 30'b000000000000000001010001100000
                ;mem[8300] <= 30'b000000000000000001010001110000
                ;mem[8301] <= 30'b000000000000000001010010000000
                ;mem[8302] <= 30'b000000000000000001010010010000
                ;mem[8303] <= 30'b000000000000000000101100100000
                ;mem[8304] <= 30'b000000000000000000101100110000
                ;mem[8305] <= 30'b000000000000000000101101000000
                ;mem[8306] <= 30'b000000000000000000101101010000
                ;mem[8307] <= 30'b000000000000000000101101100000
                ;mem[8308] <= 30'b000000000000000000101101110000
                ;mem[8309] <= 30'b000000000000000000110011100000
                ;mem[8310] <= 30'b000000000000000000110100010000
                ;mem[8311] <= 30'b000000000000000000110100100000
                ;mem[8312] <= 30'b000000000000000000110100110000
                ;mem[8313] <= 30'b000000000000000000110101000000
                ;mem[8314] <= 30'b000000000000000000110101010000
                ;mem[8315] <= 30'b000000000000000000110101100000
                ;mem[8316] <= 30'b000000000000000000111010010000
                ;mem[8317] <= 30'b000000000000000000111010100000
                ;mem[8318] <= 30'b000000001000000000000000100000
                ;mem[8319] <= 30'b000000001000000000000000110000
                ;mem[8320] <= 30'b000000001000000000000001000000
                ;mem[8321] <= 30'b000000001000000000000001010000
                ;mem[8322] <= 30'b000000001000000000000001100000
                ;mem[8323] <= 30'b000000001000000000000001110000
                ;mem[8324] <= 30'b000000001000000000000111100000
                ;mem[8325] <= 30'b000000001000000000001000010000
                ;mem[8326] <= 30'b000000001000000000001000100000
                ;mem[8327] <= 30'b000000001000000000001000110000
                ;mem[8328] <= 30'b000000001000000000001001000000
                ;mem[8329] <= 30'b000000001000000000001001010000
                ;mem[8330] <= 30'b000000001000000000001001100000
                ;mem[8331] <= 30'b000000001000000000001110010000
                ;mem[8332] <= 30'b000000001000000000001110100000
                ;mem[8333] <= 30'b000000001000000000010101010000
                ;mem[8334] <= 30'b000000001000000000010101100000
                ;mem[8335] <= 30'b000000001000000000011100010000
                ;mem[8336] <= 30'b000000001000000000100011010000
                ;mem[8337] <= 30'b000000001000000000100011100000
                ;mem[8338] <= 30'b000000001000000000101010010000
                ;mem[8339] <= 30'b000000001000000000101010100000
                ;mem[8340] <= 30'b000000001000000000101100000000
                ;mem[8341] <= 30'b000000001000000000110001010000
                ;mem[8342] <= 30'b000000001000000000110001100000
                ;mem[8343] <= 30'b000000001000000000110011000000
                ;mem[8344] <= 30'b000000001000000000110011010000
                ;mem[8345] <= 30'b000000001000000000111000100000
                ;mem[8346] <= 30'b000000001000000000111010000000
                ;mem[8347] <= 30'b000000001000000000111111100000
                ;mem[8348] <= 30'b000000001000000000111111110000
                ;mem[8349] <= 30'b000000010000000000000000000000
                ;mem[8350] <= 30'b000000010000000000000101010000
                ;mem[8351] <= 30'b000000010000000000000101100000
                ;mem[8352] <= 30'b000000010000000000000111000000
                ;mem[8353] <= 30'b000000010000000000000111010000
                ;mem[8354] <= 30'b000000010000000000001100100000
                ;mem[8355] <= 30'b000000010000000000001110000000
                ;mem[8356] <= 30'b000000010000000000010011100000
                ;mem[8357] <= 30'b000000010000000000010011110000
                ;mem[8358] <= 30'b000000010000000000010100110000
                ;mem[8359] <= 30'b000000010000000000010101000000
                ;mem[8360] <= 30'b000000010000000000011010110000
                ;mem[8361] <= 30'b000000010000000000011011000000
                ;mem[8362] <= 30'b000000010000000000011011110000
                ;mem[8363] <= 30'b000000010000000000011100000000
                ;mem[8364] <= 30'b000000010000000000100001110000
                ;mem[8365] <= 30'b000000010000000000100010000000
                ;mem[8366] <= 30'b000000010000000000100010010000
                ;mem[8367] <= 30'b000000010000000000100010100000
                ;mem[8368] <= 30'b000000010000000000100010110000
                ;mem[8369] <= 30'b000000010000000000100011000000
                ;mem[8370] <= 30'b000000010000000000101001010000
                ;mem[8371] <= 30'b000000010000000000101001110000
                ;mem[8372] <= 30'b000000010000000000101010000000
                ;mem[8373] <= 30'b000000010000000000110001000000
                ;mem[8374] <= 30'b000000010000000000111000000000
                ;mem[8375] <= 30'b000000010000000000111110110000
                ;mem[8376] <= 30'b000000010000000000111111000000
                ;mem[8377] <= 30'b000000000000000001000101000000
                ;mem[8378] <= 30'b000000000000000001001100000000
                ;mem[8379] <= 30'b000000000000000001010010110000
                ;mem[8380] <= 30'b000000000000000001010011000000
                ;mem[8381] <= 30'b000000000000000001011001110000
                ;mem[8382] <= 30'b000000000000000001011010000000
                ;mem[8383] <= 30'b000000000000000001100001000000
                ;mem[8384] <= 30'b000000000000000001101000000000
                ;mem[8385] <= 30'b000000000000000001101111000000
                ;mem[8386] <= 30'b000000000000000000011000000000
                ;mem[8387] <= 30'b000000000000000000011110110000
                ;mem[8388] <= 30'b000000000000000000011111000000
                ;mem[8389] <= 30'b000000000000000000011111010000
                ;mem[8390] <= 30'b000000000000000000011111100000
                ;mem[8391] <= 30'b000000000000000000100110000000
                ;mem[8392] <= 30'b000000000000000000100110010000
                ;mem[8393] <= 30'b000000000000000000100110100000
                ;mem[8394] <= 30'b000000000000000000100110110000
                ;mem[8395] <= 30'b000000000000000000101101010000
                ;mem[8396] <= 30'b000000000000000000101101100000
                ;mem[8397] <= 30'b000000000000000000101101110000
                ;mem[8398] <= 30'b000000000000000000101110000000
                ;mem[8399] <= 30'b000000000000000000101110010000
                ;mem[8400] <= 30'b000000000000000000110100110000
                ;mem[8401] <= 30'b000000000000000000110101000000
                ;mem[8402] <= 30'b000000000000000000110101010000
                ;mem[8403] <= 30'b000000000000000000110101100000
                ;mem[8404] <= 30'b000000000000000000111100000000
                ;mem[8405] <= 30'b000000000000000000111100010000
                ;mem[8406] <= 30'b000000000000000000111100100000
                ;mem[8407] <= 30'b000000001000000000000001010000
                ;mem[8408] <= 30'b000000001000000000000001100000
                ;mem[8409] <= 30'b000000001000000000000001110000
                ;mem[8410] <= 30'b000000001000000000000010000000
                ;mem[8411] <= 30'b000000001000000000000010010000
                ;mem[8412] <= 30'b000000001000000000001000110000
                ;mem[8413] <= 30'b000000001000000000001001000000
                ;mem[8414] <= 30'b000000001000000000001001010000
                ;mem[8415] <= 30'b000000001000000000001001100000
                ;mem[8416] <= 30'b000000001000000000010000000000
                ;mem[8417] <= 30'b000000001000000000010000010000
                ;mem[8418] <= 30'b000000001000000000010000100000
                ;mem[8419] <= 30'b000000001000000000010111010000
                ;mem[8420] <= 30'b000000001000000000010111100000
                ;mem[8421] <= 30'b000000001000000000010111110000
                ;mem[8422] <= 30'b000000001000000000011110100000
                ;mem[8423] <= 30'b000000001000000000011110110000
                ;mem[8424] <= 30'b000000001000000000100101100000
                ;mem[8425] <= 30'b000000001000000000100101110000
                ;mem[8426] <= 30'b000000001000000000101100000000
                ;mem[8427] <= 30'b000000001000000000101100010000
                ;mem[8428] <= 30'b000000001000000000101100100000
                ;mem[8429] <= 30'b000000001000000000101100110000
                ;mem[8430] <= 30'b000000001000000000110001010000
                ;mem[8431] <= 30'b000000001000000000110001100000
                ;mem[8432] <= 30'b000000001000000000110001110000
                ;mem[8433] <= 30'b000000001000000000110010000000
                ;mem[8434] <= 30'b000000001000000000110010010000
                ;mem[8435] <= 30'b000000001000000000110010110000
                ;mem[8436] <= 30'b000000001000000000110011000000
                ;mem[8437] <= 30'b000000001000000000110011010000
                ;mem[8438] <= 30'b000000001000000000110011100000
                ;mem[8439] <= 30'b000000001000000000111000010000
                ;mem[8440] <= 30'b000000001000000000111000100000
                ;mem[8441] <= 30'b000000001000000000111000110000
                ;mem[8442] <= 30'b000000001000000000111001000000
                ;mem[8443] <= 30'b000000001000000000111001010000
                ;mem[8444] <= 30'b000000001000000000111001100000
                ;mem[8445] <= 30'b000000001000000000111001110000
                ;mem[8446] <= 30'b000000001000000000111010000000
                ;mem[8447] <= 30'b000000010000000000000000000000
                ;mem[8448] <= 30'b000000010000000000000000010000
                ;mem[8449] <= 30'b000000010000000000000000100000
                ;mem[8450] <= 30'b000000010000000000000000110000
                ;mem[8451] <= 30'b000000010000000000000101010000
                ;mem[8452] <= 30'b000000010000000000000101100000
                ;mem[8453] <= 30'b000000010000000000000101110000
                ;mem[8454] <= 30'b000000010000000000000110000000
                ;mem[8455] <= 30'b000000010000000000000110010000
                ;mem[8456] <= 30'b000000010000000000000110110000
                ;mem[8457] <= 30'b000000010000000000000111000000
                ;mem[8458] <= 30'b000000010000000000000111010000
                ;mem[8459] <= 30'b000000010000000000000111100000
                ;mem[8460] <= 30'b000000010000000000001100010000
                ;mem[8461] <= 30'b000000010000000000001100100000
                ;mem[8462] <= 30'b000000010000000000001100110000
                ;mem[8463] <= 30'b000000010000000000001101000000
                ;mem[8464] <= 30'b000000010000000000001101010000
                ;mem[8465] <= 30'b000000010000000000001101100000
                ;mem[8466] <= 30'b000000010000000000001101110000
                ;mem[8467] <= 30'b000000010000000000001110000000
                ;mem[8468] <= 30'b000000010000000000010100000000
                ;mem[8469] <= 30'b000000010000000000010100010000
                ;mem[8470] <= 30'b000000010000000000010100100000
                ;mem[8471] <= 30'b000000010000000000010100110000
                ;mem[8472] <= 30'b000000010000000000010101000000
                ;mem[8473] <= 30'b000000010000000000011011100000
                ;mem[8474] <= 30'b000000010000000000011011110000
                ;mem[8475] <= 30'b000000010000000000011100000000
                ;mem[8476] <= 30'b000000010000000000100010110000
                ;mem[8477] <= 30'b000000010000000000100011000000
                ;mem[8478] <= 30'b000000010000000000101001110000
                ;mem[8479] <= 30'b000000010000000000101010000000
                ;mem[8480] <= 30'b000000010000000000101110110000
                ;mem[8481] <= 30'b000000010000000000110000010000
                ;mem[8482] <= 30'b000000010000000000110000100000
                ;mem[8483] <= 30'b000000010000000000110000110000
                ;mem[8484] <= 30'b000000010000000000110001000000
                ;mem[8485] <= 30'b000000010000000000110101100000
                ;mem[8486] <= 30'b000000010000000000110101110000
                ;mem[8487] <= 30'b000000010000000000110111000000
                ;mem[8488] <= 30'b000000010000000000110111010000
                ;mem[8489] <= 30'b000000010000000000110111100000
                ;mem[8490] <= 30'b000000010000000000110111110000
                ;mem[8491] <= 30'b000000010000000000111000000000
                ;mem[8492] <= 30'b000000010000000000111100100000
                ;mem[8493] <= 30'b000000010000000000111100110000
                ;mem[8494] <= 30'b000000010000000000111101000000
                ;mem[8495] <= 30'b000000010000000000111101010000
                ;mem[8496] <= 30'b000000010000000000111101100000
                ;mem[8497] <= 30'b000000010000000000111101110000
                ;mem[8498] <= 30'b000000010000000000111110000000
                ;mem[8499] <= 30'b000000010000000000111110010000
                ;mem[8500] <= 30'b000000000000000001000010110000
                ;mem[8501] <= 30'b000000000000000001000100010000
                ;mem[8502] <= 30'b000000000000000001000100100000
                ;mem[8503] <= 30'b000000000000000001000100110000
                ;mem[8504] <= 30'b000000000000000001000101000000
                ;mem[8505] <= 30'b000000000000000001001001100000
                ;mem[8506] <= 30'b000000000000000001001001110000
                ;mem[8507] <= 30'b000000000000000001001011000000
                ;mem[8508] <= 30'b000000000000000001001011010000
                ;mem[8509] <= 30'b000000000000000001001011100000
                ;mem[8510] <= 30'b000000000000000001001011110000
                ;mem[8511] <= 30'b000000000000000001001100000000
                ;mem[8512] <= 30'b000000000000000001010000100000
                ;mem[8513] <= 30'b000000000000000001010000110000
                ;mem[8514] <= 30'b000000000000000001010001000000
                ;mem[8515] <= 30'b000000000000000001010001010000
                ;mem[8516] <= 30'b000000000000000001010001100000
                ;mem[8517] <= 30'b000000000000000001010001110000
                ;mem[8518] <= 30'b000000000000000001010010000000
                ;mem[8519] <= 30'b000000000000000001010010010000
                ;mem[8520] <= 30'b000000000000000001010111100000
                ;mem[8521] <= 30'b000000000000000001010111110000
                ;mem[8522] <= 30'b000000000000000001011000000000
                ;mem[8523] <= 30'b000000000000000001011000010000
                ;mem[8524] <= 30'b000000000000000001011000100000
                ;mem[8525] <= 30'b000000000000000001011000110000
                ;mem[8526] <= 30'b000000000000000000110010010000
                ;mem[8527] <= 30'b000000000000000000110010100000
                ;mem[8528] <= 30'b000000000000000000110010110000
                ;mem[8529] <= 30'b000000000000000000110011000000
                ;mem[8530] <= 30'b000000000000000000110011010000
                ;mem[8531] <= 30'b000000000000000000110011100000
                ;mem[8532] <= 30'b000000000000000000110011110000
                ;mem[8533] <= 30'b000000000000000000110100000000
                ;mem[8534] <= 30'b000000000000000000110100010000
                ;mem[8535] <= 30'b000000000000000000110100100000
                ;mem[8536] <= 30'b000000000000000000110101010000
                ;mem[8537] <= 30'b000000000000000000111001010000
                ;mem[8538] <= 30'b000000000000000000111001100000
                ;mem[8539] <= 30'b000000000000000000111001110000
                ;mem[8540] <= 30'b000000000000000000111010000000
                ;mem[8541] <= 30'b000000000000000000111010010000
                ;mem[8542] <= 30'b000000000000000000111010100000
                ;mem[8543] <= 30'b000000000000000000111010110000
                ;mem[8544] <= 30'b000000000000000000111011000000
                ;mem[8545] <= 30'b000000000000000000111011010000
                ;mem[8546] <= 30'b000000000000000000111011100000
                ;mem[8547] <= 30'b000000000000000000111011110000
                ;mem[8548] <= 30'b000000000000000000111100000000
                ;mem[8549] <= 30'b000000000000000000111100010000
                ;mem[8550] <= 30'b000000000000000000111100100000
                ;mem[8551] <= 30'b000000000000000000111100110000
                ;mem[8552] <= 30'b000000000000000000111101000000
                ;mem[8553] <= 30'b000000000000000000111101010000
                ;mem[8554] <= 30'b000000000000000000111101100000
                ;mem[8555] <= 30'b000000001000000000000110010000
                ;mem[8556] <= 30'b000000001000000000000110100000
                ;mem[8557] <= 30'b000000001000000000000110110000
                ;mem[8558] <= 30'b000000001000000000000111000000
                ;mem[8559] <= 30'b000000001000000000000111010000
                ;mem[8560] <= 30'b000000001000000000000111100000
                ;mem[8561] <= 30'b000000001000000000000111110000
                ;mem[8562] <= 30'b000000001000000000001000000000
                ;mem[8563] <= 30'b000000001000000000001000010000
                ;mem[8564] <= 30'b000000001000000000001000100000
                ;mem[8565] <= 30'b000000001000000000001001010000
                ;mem[8566] <= 30'b000000001000000000001101010000
                ;mem[8567] <= 30'b000000001000000000001101100000
                ;mem[8568] <= 30'b000000001000000000001101110000
                ;mem[8569] <= 30'b000000001000000000001110000000
                ;mem[8570] <= 30'b000000001000000000001110010000
                ;mem[8571] <= 30'b000000001000000000001110100000
                ;mem[8572] <= 30'b000000001000000000001110110000
                ;mem[8573] <= 30'b000000001000000000001111000000
                ;mem[8574] <= 30'b000000001000000000001111010000
                ;mem[8575] <= 30'b000000001000000000001111100000
                ;mem[8576] <= 30'b000000001000000000001111110000
                ;mem[8577] <= 30'b000000001000000000010000000000
                ;mem[8578] <= 30'b000000001000000000010000010000
                ;mem[8579] <= 30'b000000001000000000010000100000
                ;mem[8580] <= 30'b000000001000000000010000110000
                ;mem[8581] <= 30'b000000001000000000010001000000
                ;mem[8582] <= 30'b000000001000000000010001010000
                ;mem[8583] <= 30'b000000001000000000010001100000
                ;mem[8584] <= 30'b000000001000000000010110000000
                ;mem[8585] <= 30'b000000001000000000010110010000
                ;mem[8586] <= 30'b000000001000000000010110100000
                ;mem[8587] <= 30'b000000001000000000010110110000
                ;mem[8588] <= 30'b000000001000000000010111000000
                ;mem[8589] <= 30'b000000001000000000010111010000
                ;mem[8590] <= 30'b000000001000000000010111100000
                ;mem[8591] <= 30'b000000001000000000010111110000
                ;mem[8592] <= 30'b000000001000000000011000000000
                ;mem[8593] <= 30'b000000001000000000011000010000
                ;mem[8594] <= 30'b000000001000000000011000100000
                ;mem[8595] <= 30'b000000001000000000011110110000
                ;mem[8596] <= 30'b000000001000000000011111000000
                ;mem[8597] <= 30'b000000001000000000011111010000
                ;mem[8598] <= 30'b000000001000000000011111100000
                ;mem[8599] <= 30'b000000001000000000100101110000
                ;mem[8600] <= 30'b000000001000000000100110000000
                ;mem[8601] <= 30'b000000001000000000100110010000
                ;mem[8602] <= 30'b000000001000000000101100100000
                ;mem[8603] <= 30'b000000001000000000101100110000
                ;mem[8604] <= 30'b000000001000000000101101000000
                ;mem[8605] <= 30'b000000001000000000110011010000
                ;mem[8606] <= 30'b000000001000000000110011100000
                ;mem[8607] <= 30'b000000001000000000110011110000
                ;mem[8608] <= 30'b000000001000000000111000010000
                ;mem[8609] <= 30'b000000001000000000111000100000
                ;mem[8610] <= 30'b000000001000000000111000110000
                ;mem[8611] <= 30'b000000001000000000111001000000
                ;mem[8612] <= 30'b000000001000000000111001010000
                ;mem[8613] <= 30'b000000001000000000111001100000
                ;mem[8614] <= 30'b000000001000000000111001110000
                ;mem[8615] <= 30'b000000001000000000111010000000
                ;mem[8616] <= 30'b000000001000000000111010010000
                ;mem[8617] <= 30'b000000001000000000111010100000
                ;mem[8618] <= 30'b000000001000000000111010110000
                ;mem[8619] <= 30'b000000001000000000111111010000
                ;mem[8620] <= 30'b000000001000000000111111100000
                ;mem[8621] <= 30'b000000001000000000111111110000
                ;mem[8622] <= 30'b000000010000000000000000100000
                ;mem[8623] <= 30'b000000010000000000000000110000
                ;mem[8624] <= 30'b000000010000000000000001000000
                ;mem[8625] <= 30'b000000010000000000000111010000
                ;mem[8626] <= 30'b000000010000000000000111100000
                ;mem[8627] <= 30'b000000010000000000000111110000
                ;mem[8628] <= 30'b000000010000000000001100010000
                ;mem[8629] <= 30'b000000010000000000001100100000
                ;mem[8630] <= 30'b000000010000000000001100110000
                ;mem[8631] <= 30'b000000010000000000001101000000
                ;mem[8632] <= 30'b000000010000000000001101010000
                ;mem[8633] <= 30'b000000010000000000001101100000
                ;mem[8634] <= 30'b000000010000000000001101110000
                ;mem[8635] <= 30'b000000010000000000001110000000
                ;mem[8636] <= 30'b000000010000000000001110010000
                ;mem[8637] <= 30'b000000010000000000001110100000
                ;mem[8638] <= 30'b000000010000000000001110110000
                ;mem[8639] <= 30'b000000010000000000010011010000
                ;mem[8640] <= 30'b000000010000000000010011100000
                ;mem[8641] <= 30'b000000010000000000010011110000
                ;mem[8642] <= 30'b000000010000000000010100000000
                ;mem[8643] <= 30'b000000010000000000010100010000
                ;mem[8644] <= 30'b000000010000000000010100100000
                ;mem[8645] <= 30'b000000010000000000010100110000
                ;mem[8646] <= 30'b000000010000000000010101000000
                ;mem[8647] <= 30'b000000010000000000010101010000
                ;mem[8648] <= 30'b000000010000000000010101100000
                ;mem[8649] <= 30'b000000010000000000010101110000
                ;mem[8650] <= 30'b000000010000000000010110000000
                ;mem[8651] <= 30'b000000010000000000010110010000
                ;mem[8652] <= 30'b000000010000000000010110100000
                ;mem[8653] <= 30'b000000010000000000011010110000
                ;mem[8654] <= 30'b000000010000000000011011000000
                ;mem[8655] <= 30'b000000010000000000011011010000
                ;mem[8656] <= 30'b000000010000000000011011100000
                ;mem[8657] <= 30'b000000010000000000011011110000
                ;mem[8658] <= 30'b000000010000000000011100000000
                ;mem[8659] <= 30'b000000010000000000011100010000
                ;mem[8660] <= 30'b000000010000000000011100100000
                ;mem[8661] <= 30'b000000010000000000011100110000
                ;mem[8662] <= 30'b000000010000000000011101000000
                ;mem[8663] <= 30'b000000010000000000011101010000
                ;mem[8664] <= 30'b000000010000000000011101100000
                ;mem[8665] <= 30'b000000010000000000100010010000
                ;mem[8666] <= 30'b000000010000000000100010100000
                ;mem[8667] <= 30'b000000010000000000100010110000
                ;mem[8668] <= 30'b000000010000000000100011000000
                ;mem[8669] <= 30'b000000010000000000100011010000
                ;mem[8670] <= 30'b000000010000000000101001000000
                ;mem[8671] <= 30'b000000010000000000101001010000
                ;mem[8672] <= 30'b000000010000000000101001100000
                ;mem[8673] <= 30'b000000010000000000101001110000
                ;mem[8674] <= 30'b000000010000000000101111110000
                ;mem[8675] <= 30'b000000010000000000110000000000
                ;mem[8676] <= 30'b000000010000000000110000010000
                ;mem[8677] <= 30'b000000010000000000110110110000
                ;mem[8678] <= 30'b000000010000000000110111000000
                ;mem[8679] <= 30'b000000010000000000110111010000
                ;mem[8680] <= 30'b000000010000000000111101100000
                ;mem[8681] <= 30'b000000010000000000111101110000
                ;mem[8682] <= 30'b000000010000000000111110000000
                ;mem[8683] <= 30'b000000000000000001000011110000
                ;mem[8684] <= 30'b000000000000000001000100000000
                ;mem[8685] <= 30'b000000000000000001000100010000
                ;mem[8686] <= 30'b000000000000000001001010110000
                ;mem[8687] <= 30'b000000000000000001001011000000
                ;mem[8688] <= 30'b000000000000000001001011010000
                ;mem[8689] <= 30'b000000000000000001010001100000
                ;mem[8690] <= 30'b000000000000000001010001110000
                ;mem[8691] <= 30'b000000000000000001010010000000
                ;mem[8692] <= 30'b000000000000000001011000100000
                ;mem[8693] <= 30'b000000000000000001011000110000
                ;mem[8694] <= 30'b000000000000000001011111010000
                ;mem[8695] <= 30'b000000000000000001011111100000
                ;mem[8696] <= 30'b000000000000000001100110000000
                ;mem[8697] <= 30'b000000000000000001100110010000
                ;mem[8698] <= 30'b000000000000000001100110100000
                ;mem[8699] <= 30'b000000000000000001101100110000
                ;mem[8700] <= 30'b000000000000000001101101000000
                ;mem[8701] <= 30'b000000000000000001101101010000
                ;mem[8702] <= 30'b000000000000000001110011110000
                ;mem[8703] <= 30'b000000000000000001110100000000
                ;mem[8704] <= 30'b000000000000000001110100010000
                ;mem[8705] <= 30'b000000000000000000100111000000
                ;mem[8706] <= 30'b000000000000000000101110000000
                ;mem[8707] <= 30'b000000000000000000101110010000
                ;mem[8708] <= 30'b000000000000000000110101000000
                ;mem[8709] <= 30'b000000000000000000110101010000
                ;mem[8710] <= 30'b000000000000000000111011000000
                ;mem[8711] <= 30'b000000000000000000111100000000
                ;mem[8712] <= 30'b000000000000000000111100010000
                ;mem[8713] <= 30'b000000001000000000000010000000
                ;mem[8714] <= 30'b000000001000000000000010010000
                ;mem[8715] <= 30'b000000001000000000001001000000
                ;mem[8716] <= 30'b000000001000000000001001010000
                ;mem[8717] <= 30'b000000001000000000001111000000
                ;mem[8718] <= 30'b000000001000000000010000000000
                ;mem[8719] <= 30'b000000001000000000010000010000
                ;mem[8720] <= 30'b000000001000000000010110000000
                ;mem[8721] <= 30'b000000001000000000010111000000
                ;mem[8722] <= 30'b000000001000000000010111010000
                ;mem[8723] <= 30'b000000001000000000011101000000
                ;mem[8724] <= 30'b000000001000000000011110000000
                ;mem[8725] <= 30'b000000001000000000011110010000
                ;mem[8726] <= 30'b000000001000000000100011110000
                ;mem[8727] <= 30'b000000001000000000100100000000
                ;mem[8728] <= 30'b000000001000000000100101000000
                ;mem[8729] <= 30'b000000001000000000100101010000
                ;mem[8730] <= 30'b000000001000000000101010110000
                ;mem[8731] <= 30'b000000001000000000101011000000
                ;mem[8732] <= 30'b000000001000000000101100000000
                ;mem[8733] <= 30'b000000001000000000101100010000
                ;mem[8734] <= 30'b000000001000000000110001100000
                ;mem[8735] <= 30'b000000001000000000110001110000
                ;mem[8736] <= 30'b000000001000000000110010000000
                ;mem[8737] <= 30'b000000001000000000110010010000
                ;mem[8738] <= 30'b000000001000000000110011000000
                ;mem[8739] <= 30'b000000001000000000110011010000
                ;mem[8740] <= 30'b000000001000000000111000100000
                ;mem[8741] <= 30'b000000001000000000111000110000
                ;mem[8742] <= 30'b000000001000000000111001000000
                ;mem[8743] <= 30'b000000001000000000111001010000
                ;mem[8744] <= 30'b000000001000000000111001100000
                ;mem[8745] <= 30'b000000001000000000111001110000
                ;mem[8746] <= 30'b000000001000000000111010000000
                ;mem[8747] <= 30'b000000001000000000111010010000
                ;mem[8748] <= 30'b000000001000000000111111100000
                ;mem[8749] <= 30'b000000001000000000111111110000
                ;mem[8750] <= 30'b000000010000000000000000000000
                ;mem[8751] <= 30'b000000010000000000000000010000
                ;mem[8752] <= 30'b000000010000000000000101100000
                ;mem[8753] <= 30'b000000010000000000000101110000
                ;mem[8754] <= 30'b000000010000000000000110000000
                ;mem[8755] <= 30'b000000010000000000000110010000
                ;mem[8756] <= 30'b000000010000000000000111000000
                ;mem[8757] <= 30'b000000010000000000000111010000
                ;mem[8758] <= 30'b000000010000000000001100100000
                ;mem[8759] <= 30'b000000010000000000001100110000
                ;mem[8760] <= 30'b000000010000000000001101000000
                ;mem[8761] <= 30'b000000010000000000001101010000
                ;mem[8762] <= 30'b000000010000000000001101100000
                ;mem[8763] <= 30'b000000010000000000001101110000
                ;mem[8764] <= 30'b000000010000000000001110000000
                ;mem[8765] <= 30'b000000010000000000001110010000
                ;mem[8766] <= 30'b000000010000000000010011100000
                ;mem[8767] <= 30'b000000010000000000010011110000
                ;mem[8768] <= 30'b000000010000000000010100000000
                ;mem[8769] <= 30'b000000010000000000010101000000
                ;mem[8770] <= 30'b000000010000000000010101010000
                ;mem[8771] <= 30'b000000010000000000011010100000
                ;mem[8772] <= 30'b000000010000000000011100000000
                ;mem[8773] <= 30'b000000010000000000011100010000
                ;mem[8774] <= 30'b000000010000000000100011000000
                ;mem[8775] <= 30'b000000010000000000100011010000
                ;mem[8776] <= 30'b000000010000000000101010000000
                ;mem[8777] <= 30'b000000010000000000101010010000
                ;mem[8778] <= 30'b000000010000000000110001000000
                ;mem[8779] <= 30'b000000010000000000110001010000
                ;mem[8780] <= 30'b000000010000000000111000000000
                ;mem[8781] <= 30'b000000010000000000111110110000
                ;mem[8782] <= 30'b000000010000000000111111000000
                ;mem[8783] <= 30'b000000000000000001000101000000
                ;mem[8784] <= 30'b000000000000000001000101010000
                ;mem[8785] <= 30'b000000000000000001001100000000
                ;mem[8786] <= 30'b000000000000000001010010110000
                ;mem[8787] <= 30'b000000000000000001010011000000
                ;mem[8788] <= 30'b000000000000000001011001110000
                ;mem[8789] <= 30'b000000000000000001011010000000
                ;mem[8790] <= 30'b000000000000000001100000110000
                ;mem[8791] <= 30'b000000000000000001100001000000
                ;mem[8792] <= 30'b000000000000000000010001010000
                ;mem[8793] <= 30'b000000000000000000011000000000
                ;mem[8794] <= 30'b000000000000000000011000010000
                ;mem[8795] <= 30'b000000000000000000011110110000
                ;mem[8796] <= 30'b000000000000000000011111000000
                ;mem[8797] <= 30'b000000000000000000011111010000
                ;mem[8798] <= 30'b000000000000000000100101100000
                ;mem[8799] <= 30'b000000000000000000100101110000
                ;mem[8800] <= 30'b000000000000000000100110000000
                ;mem[8801] <= 30'b000000000000000000101100100000
                ;mem[8802] <= 30'b000000000000000000110011010000
                ;mem[8803] <= 30'b000000000000000000110011100000
                ;mem[8804] <= 30'b000000000000000000111010010000
                ;mem[8805] <= 30'b000000000000000000111100110000
                ;mem[8806] <= 30'b000000000000000000111101000000
                ;mem[8807] <= 30'b000000000000000000111101010000
                ;mem[8808] <= 30'b000000001000000000000000100000
                ;mem[8809] <= 30'b000000001000000000000111010000
                ;mem[8810] <= 30'b000000001000000000000111100000
                ;mem[8811] <= 30'b000000001000000000001110010000
                ;mem[8812] <= 30'b000000001000000000010000110000
                ;mem[8813] <= 30'b000000001000000000010001000000
                ;mem[8814] <= 30'b000000001000000000010001010000
                ;mem[8815] <= 30'b000000001000000000010101000000
                ;mem[8816] <= 30'b000000001000000000010101010000
                ;mem[8817] <= 30'b000000001000000000010111010000
                ;mem[8818] <= 30'b000000001000000000010111100000
                ;mem[8819] <= 30'b000000001000000000010111110000
                ;mem[8820] <= 30'b000000001000000000011000000000
                ;mem[8821] <= 30'b000000001000000000011000010000
                ;mem[8822] <= 30'b000000001000000000011100000000
                ;mem[8823] <= 30'b000000001000000000011100010000
                ;mem[8824] <= 30'b000000001000000000011110000000
                ;mem[8825] <= 30'b000000001000000000011110010000
                ;mem[8826] <= 30'b000000001000000000011110100000
                ;mem[8827] <= 30'b000000001000000000011111000000
                ;mem[8828] <= 30'b000000001000000000011111010000
                ;mem[8829] <= 30'b000000001000000000100011000000
                ;mem[8830] <= 30'b000000001000000000100100110000
                ;mem[8831] <= 30'b000000001000000000100101000000
                ;mem[8832] <= 30'b000000001000000000100101010000
                ;mem[8833] <= 30'b000000001000000000100110000000
                ;mem[8834] <= 30'b000000001000000000100110010000
                ;mem[8835] <= 30'b000000001000000000101001110000
                ;mem[8836] <= 30'b000000001000000000101010000000
                ;mem[8837] <= 30'b000000001000000000101011110000
                ;mem[8838] <= 30'b000000001000000000101100000000
                ;mem[8839] <= 30'b000000001000000000101101000000
                ;mem[8840] <= 30'b000000001000000000101101010000
                ;mem[8841] <= 30'b000000001000000000110000110000
                ;mem[8842] <= 30'b000000001000000000110001000000
                ;mem[8843] <= 30'b000000001000000000110010100000
                ;mem[8844] <= 30'b000000001000000000110010110000
                ;mem[8845] <= 30'b000000001000000000110100000000
                ;mem[8846] <= 30'b000000001000000000110100010000
                ;mem[8847] <= 30'b000000001000000000110111110000
                ;mem[8848] <= 30'b000000001000000000111000000000
                ;mem[8849] <= 30'b000000001000000000111001100000
                ;mem[8850] <= 30'b000000001000000000111001110000
                ;mem[8851] <= 30'b000000001000000000111011000000
                ;mem[8852] <= 30'b000000001000000000111011010000
                ;mem[8853] <= 30'b000000001000000000111110110000
                ;mem[8854] <= 30'b000000010000000000000000000000
                ;mem[8855] <= 30'b000000010000000000000001000000
                ;mem[8856] <= 30'b000000010000000000000001010000
                ;mem[8857] <= 30'b000000010000000000000100110000
                ;mem[8858] <= 30'b000000010000000000000101000000
                ;mem[8859] <= 30'b000000010000000000000110100000
                ;mem[8860] <= 30'b000000010000000000000110110000
                ;mem[8861] <= 30'b000000010000000000001000000000
                ;mem[8862] <= 30'b000000010000000000001000010000
                ;mem[8863] <= 30'b000000010000000000001011110000
                ;mem[8864] <= 30'b000000010000000000001100000000
                ;mem[8865] <= 30'b000000010000000000001101100000
                ;mem[8866] <= 30'b000000010000000000001101110000
                ;mem[8867] <= 30'b000000010000000000001111000000
                ;mem[8868] <= 30'b000000010000000000001111010000
                ;mem[8869] <= 30'b000000010000000000010010110000
                ;mem[8870] <= 30'b000000010000000000010100100000
                ;mem[8871] <= 30'b000000010000000000010100110000
                ;mem[8872] <= 30'b000000010000000000010101110000
                ;mem[8873] <= 30'b000000010000000000010110000000
                ;mem[8874] <= 30'b000000010000000000011001110000
                ;mem[8875] <= 30'b000000010000000000011010000000
                ;mem[8876] <= 30'b000000010000000000011011100000
                ;mem[8877] <= 30'b000000010000000000011100110000
                ;mem[8878] <= 30'b000000010000000000011101000000
                ;mem[8879] <= 30'b000000010000000000100000110000
                ;mem[8880] <= 30'b000000010000000000100001000000
                ;mem[8881] <= 30'b000000010000000000100010100000
                ;mem[8882] <= 30'b000000010000000000100011100000
                ;mem[8883] <= 30'b000000010000000000100011110000
                ;mem[8884] <= 30'b000000010000000000101000000000
                ;mem[8885] <= 30'b000000010000000000101000010000
                ;mem[8886] <= 30'b000000010000000000101001100000
                ;mem[8887] <= 30'b000000010000000000101001110000
                ;mem[8888] <= 30'b000000010000000000101010010000
                ;mem[8889] <= 30'b000000010000000000101010100000
                ;mem[8890] <= 30'b000000010000000000101111000000
                ;mem[8891] <= 30'b000000010000000000101111010000
                ;mem[8892] <= 30'b000000010000000000101111100000
                ;mem[8893] <= 30'b000000010000000000110000100000
                ;mem[8894] <= 30'b000000010000000000110000110000
                ;mem[8895] <= 30'b000000010000000000110001000000
                ;mem[8896] <= 30'b000000010000000000110001010000
                ;mem[8897] <= 30'b000000010000000000110110010000
                ;mem[8898] <= 30'b000000010000000000110110100000
                ;mem[8899] <= 30'b000000010000000000110110110000
                ;mem[8900] <= 30'b000000010000000000110111000000
                ;mem[8901] <= 30'b000000010000000000110111010000
                ;mem[8902] <= 30'b000000010000000000110111100000
                ;mem[8903] <= 30'b000000010000000000110111110000
                ;mem[8904] <= 30'b000000010000000000111000000000
                ;mem[8905] <= 30'b000000010000000000111000010000
                ;mem[8906] <= 30'b000000010000000000111101100000
                ;mem[8907] <= 30'b000000010000000000111101110000
                ;mem[8908] <= 30'b000000010000000000111110000000
                ;mem[8909] <= 30'b000000010000000000111110010000
                ;mem[8910] <= 30'b000000010000000000111110100000
                ;mem[8911] <= 30'b000000010000000000111110110000
                ;mem[8912] <= 30'b000000010000000000111111000000
                ;mem[8913] <= 30'b000000000000000001000011000000
                ;mem[8914] <= 30'b000000000000000001000011010000
                ;mem[8915] <= 30'b000000000000000001000011100000
                ;mem[8916] <= 30'b000000000000000001000100100000
                ;mem[8917] <= 30'b000000000000000001000100110000
                ;mem[8918] <= 30'b000000000000000001000101000000
                ;mem[8919] <= 30'b000000000000000001000101010000
                ;mem[8920] <= 30'b000000000000000001001010010000
                ;mem[8921] <= 30'b000000000000000001001010100000
                ;mem[8922] <= 30'b000000000000000001001010110000
                ;mem[8923] <= 30'b000000000000000001001011000000
                ;mem[8924] <= 30'b000000000000000001001011010000
                ;mem[8925] <= 30'b000000000000000001001011100000
                ;mem[8926] <= 30'b000000000000000001001011110000
                ;mem[8927] <= 30'b000000000000000001001100000000
                ;mem[8928] <= 30'b000000000000000001001100010000
                ;mem[8929] <= 30'b000000000000000001010001100000
                ;mem[8930] <= 30'b000000000000000001010001110000
                ;mem[8931] <= 30'b000000000000000001010010000000
                ;mem[8932] <= 30'b000000000000000001010010010000
                ;mem[8933] <= 30'b000000000000000001010010100000
                ;mem[8934] <= 30'b000000000000000001010010110000
                ;mem[8935] <= 30'b000000000000000001010011000000
                ;mem[8936] <= 30'b000000000000000000101000010000
                ;mem[8937] <= 30'b000000000000000000101000100000
                ;mem[8938] <= 30'b000000000000000000101111000000
                ;mem[8939] <= 30'b000000000000000000101111010000
                ;mem[8940] <= 30'b000000000000000000101111100000
                ;mem[8941] <= 30'b000000000000000000110101110000
                ;mem[8942] <= 30'b000000000000000000110110000000
                ;mem[8943] <= 30'b000000000000000000110110010000
                ;mem[8944] <= 30'b000000000000000000111100100000
                ;mem[8945] <= 30'b000000000000000000111100110000
                ;mem[8946] <= 30'b000000000000000000111101000000
                ;mem[8947] <= 30'b000000001000000000000011000000
                ;mem[8948] <= 30'b000000001000000000000011010000
                ;mem[8949] <= 30'b000000001000000000000011100000
                ;mem[8950] <= 30'b000000001000000000001001110000
                ;mem[8951] <= 30'b000000001000000000001010000000
                ;mem[8952] <= 30'b000000001000000000001010010000
                ;mem[8953] <= 30'b000000001000000000010000100000
                ;mem[8954] <= 30'b000000001000000000010000110000
                ;mem[8955] <= 30'b000000001000000000010001000000
                ;mem[8956] <= 30'b000000001000000000010101000000
                ;mem[8957] <= 30'b000000001000000000010101010000
                ;mem[8958] <= 30'b000000001000000000010111110000
                ;mem[8959] <= 30'b000000001000000000011000000000
                ;mem[8960] <= 30'b000000001000000000011011110000
                ;mem[8961] <= 30'b000000001000000000011100000000
                ;mem[8962] <= 30'b000000001000000000011110100000
                ;mem[8963] <= 30'b000000001000000000011110110000
                ;mem[8964] <= 30'b000000001000000000100010010000
                ;mem[8965] <= 30'b000000001000000000100010100000
                ;mem[8966] <= 30'b000000001000000000100010110000
                ;mem[8967] <= 30'b000000001000000000100101010000
                ;mem[8968] <= 30'b000000001000000000100101100000
                ;mem[8969] <= 30'b000000001000000000100101110000
                ;mem[8970] <= 30'b000000001000000000101001010000
                ;mem[8971] <= 30'b000000001000000000101001100000
                ;mem[8972] <= 30'b000000001000000000101100010000
                ;mem[8973] <= 30'b000000001000000000101100100000
                ;mem[8974] <= 30'b000000001000000000101100110000
                ;mem[8975] <= 30'b000000001000000000110000010000
                ;mem[8976] <= 30'b000000001000000000110000100000
                ;mem[8977] <= 30'b000000001000000000110011010000
                ;mem[8978] <= 30'b000000001000000000110011100000
                ;mem[8979] <= 30'b000000001000000000110111010000
                ;mem[8980] <= 30'b000000001000000000110111100000
                ;mem[8981] <= 30'b000000001000000000110111110000
                ;mem[8982] <= 30'b000000001000000000111010010000
                ;mem[8983] <= 30'b000000001000000000111010100000
                ;mem[8984] <= 30'b000000001000000000111110010000
                ;mem[8985] <= 30'b000000001000000000111110100000
                ;mem[8986] <= 30'b000000001000000000111110110000
                ;mem[8987] <= 30'b000000001000000000111111000000
                ;mem[8988] <= 30'b000000010000000000000000010000
                ;mem[8989] <= 30'b000000010000000000000000100000
                ;mem[8990] <= 30'b000000010000000000000000110000
                ;mem[8991] <= 30'b000000010000000000000100010000
                ;mem[8992] <= 30'b000000010000000000000100100000
                ;mem[8993] <= 30'b000000010000000000000111010000
                ;mem[8994] <= 30'b000000010000000000000111100000
                ;mem[8995] <= 30'b000000010000000000001011010000
                ;mem[8996] <= 30'b000000010000000000001011100000
                ;mem[8997] <= 30'b000000010000000000001011110000
                ;mem[8998] <= 30'b000000010000000000001110010000
                ;mem[8999] <= 30'b000000010000000000001110100000
                ;mem[9000] <= 30'b000000010000000000010010010000
                ;mem[9001] <= 30'b000000010000000000010010100000
                ;mem[9002] <= 30'b000000010000000000010010110000
                ;mem[9003] <= 30'b000000010000000000010011000000
                ;mem[9004] <= 30'b000000010000000000010100110000
                ;mem[9005] <= 30'b000000010000000000010101000000
                ;mem[9006] <= 30'b000000010000000000010101010000
                ;mem[9007] <= 30'b000000010000000000010101100000
                ;mem[9008] <= 30'b000000010000000000011001100000
                ;mem[9009] <= 30'b000000010000000000011001110000
                ;mem[9010] <= 30'b000000010000000000011010000000
                ;mem[9011] <= 30'b000000010000000000011010010000
                ;mem[9012] <= 30'b000000010000000000011010100000
                ;mem[9013] <= 30'b000000010000000000011010110000
                ;mem[9014] <= 30'b000000010000000000011011000000
                ;mem[9015] <= 30'b000000010000000000011011010000
                ;mem[9016] <= 30'b000000010000000000011011100000
                ;mem[9017] <= 30'b000000010000000000011011110000
                ;mem[9018] <= 30'b000000010000000000011100000000
                ;mem[9019] <= 30'b000000010000000000011100010000
                ;mem[9020] <= 30'b000000010000000000011100100000
                ;mem[9021] <= 30'b000000010000000000100000110000
                ;mem[9022] <= 30'b000000010000000000100001000000
                ;mem[9023] <= 30'b000000010000000000100001010000
                ;mem[9024] <= 30'b000000010000000000100001100000
                ;mem[9025] <= 30'b000000010000000000100001110000
                ;mem[9026] <= 30'b000000010000000000100010000000
                ;mem[9027] <= 30'b000000010000000000100010010000
                ;mem[9028] <= 30'b000000010000000000100010100000
                ;mem[9029] <= 30'b000000010000000000100010110000
                ;mem[9030] <= 30'b000000010000000000100011000000
                ;mem[9031] <= 30'b000000010000000000100011010000
                ;mem[9032] <= 30'b000000010000000000101000010000
                ;mem[9033] <= 30'b000000010000000000101010000000
                ;mem[9034] <= 30'b000000010000000000101010010000
                ;mem[9035] <= 30'b000000010000000000110001000000
                ;mem[9036] <= 30'b000000010000000000110001010000
                ;mem[9037] <= 30'b000000010000000000110111110000
                ;mem[9038] <= 30'b000000010000000000111000000000
                ;mem[9039] <= 30'b000000010000000000111000010000
                ;mem[9040] <= 30'b000000010000000000111110110000
                ;mem[9041] <= 30'b000000010000000000111111000000
                ;mem[9042] <= 30'b000000010000000000111111010000
                ;mem[9043] <= 30'b000000000000000001000101000000
                ;mem[9044] <= 30'b000000000000000001000101010000
                ;mem[9045] <= 30'b000000000000000001001011110000
                ;mem[9046] <= 30'b000000000000000001001100000000
                ;mem[9047] <= 30'b000000000000000001001100010000
                ;mem[9048] <= 30'b000000000000000001010010110000
                ;mem[9049] <= 30'b000000000000000001010011000000
                ;mem[9050] <= 30'b000000000000000001010011010000
                ;mem[9051] <= 30'b000000000000000001011001110000
                ;mem[9052] <= 30'b000000000000000001011010000000
                ;mem[9053] <= 30'b000000000000000001011010010000
                ;mem[9054] <= 30'b000000000000000001100000110000
                ;mem[9055] <= 30'b000000000000000001100001000000
                ;mem[9056] <= 30'b000000000000000001100111110000
                ;mem[9057] <= 30'b000000000000000000100101010000
                ;mem[9058] <= 30'b000000000000000000100101100000
                ;mem[9059] <= 30'b000000000000000000100101110000
                ;mem[9060] <= 30'b000000000000000000100110000000
                ;mem[9061] <= 30'b000000000000000000100110010000
                ;mem[9062] <= 30'b000000000000000000100110100000
                ;mem[9063] <= 30'b000000000000000000100110110000
                ;mem[9064] <= 30'b000000000000000000100111000000
                ;mem[9065] <= 30'b000000000000000000101100000000
                ;mem[9066] <= 30'b000000000000000000101100010000
                ;mem[9067] <= 30'b000000000000000000101100100000
                ;mem[9068] <= 30'b000000000000000000101100110000
                ;mem[9069] <= 30'b000000000000000000101101000000
                ;mem[9070] <= 30'b000000000000000000101101010000
                ;mem[9071] <= 30'b000000000000000000101101100000
                ;mem[9072] <= 30'b000000000000000000101101110000
                ;mem[9073] <= 30'b000000000000000000101110000000
                ;mem[9074] <= 30'b000000000000000000101110010000
                ;mem[9075] <= 30'b000000000000000000110010110000
                ;mem[9076] <= 30'b000000000000000000110011000000
                ;mem[9077] <= 30'b000000000000000000110011010000
                ;mem[9078] <= 30'b000000000000000000110011100000
                ;mem[9079] <= 30'b000000000000000000110011110000
                ;mem[9080] <= 30'b000000000000000000110100000000
                ;mem[9081] <= 30'b000000000000000000110100010000
                ;mem[9082] <= 30'b000000000000000000110100100000
                ;mem[9083] <= 30'b000000000000000000110100110000
                ;mem[9084] <= 30'b000000000000000000110101000000
                ;mem[9085] <= 30'b000000000000000000110101010000
                ;mem[9086] <= 30'b000000000000000000110101100000
                ;mem[9087] <= 30'b000000000000000000111010000000
                ;mem[9088] <= 30'b000000000000000000111010010000
                ;mem[9089] <= 30'b000000000000000000111010100000
                ;mem[9090] <= 30'b000000000000000000111010110000
                ;mem[9091] <= 30'b000000000000000000111011100000
                ;mem[9092] <= 30'b000000000000000000111011110000
                ;mem[9093] <= 30'b000000000000000000111100000000
                ;mem[9094] <= 30'b000000000000000000111100010000
                ;mem[9095] <= 30'b000000000000000000111100100000
                ;mem[9096] <= 30'b000000000000000000111100110000
                ;mem[9097] <= 30'b000000001000000000000000000000
                ;mem[9098] <= 30'b000000001000000000000000010000
                ;mem[9099] <= 30'b000000001000000000000000100000
                ;mem[9100] <= 30'b000000001000000000000000110000
                ;mem[9101] <= 30'b000000001000000000000001000000
                ;mem[9102] <= 30'b000000001000000000000001010000
                ;mem[9103] <= 30'b000000001000000000000001100000
                ;mem[9104] <= 30'b000000001000000000000001110000
                ;mem[9105] <= 30'b000000001000000000000010000000
                ;mem[9106] <= 30'b000000001000000000000010010000
                ;mem[9107] <= 30'b000000001000000000000110110000
                ;mem[9108] <= 30'b000000001000000000000111000000
                ;mem[9109] <= 30'b000000001000000000000111010000
                ;mem[9110] <= 30'b000000001000000000000111100000
                ;mem[9111] <= 30'b000000001000000000000111110000
                ;mem[9112] <= 30'b000000001000000000001000000000
                ;mem[9113] <= 30'b000000001000000000001000010000
                ;mem[9114] <= 30'b000000001000000000001000100000
                ;mem[9115] <= 30'b000000001000000000001000110000
                ;mem[9116] <= 30'b000000001000000000001001000000
                ;mem[9117] <= 30'b000000001000000000001001010000
                ;mem[9118] <= 30'b000000001000000000001001100000
                ;mem[9119] <= 30'b000000001000000000001110000000
                ;mem[9120] <= 30'b000000001000000000001110010000
                ;mem[9121] <= 30'b000000001000000000001110100000
                ;mem[9122] <= 30'b000000001000000000001110110000
                ;mem[9123] <= 30'b000000001000000000001111100000
                ;mem[9124] <= 30'b000000001000000000001111110000
                ;mem[9125] <= 30'b000000001000000000010000000000
                ;mem[9126] <= 30'b000000001000000000010000010000
                ;mem[9127] <= 30'b000000001000000000010000100000
                ;mem[9128] <= 30'b000000001000000000010000110000
                ;mem[9129] <= 30'b000000001000000000010110110000
                ;mem[9130] <= 30'b000000001000000000010111000000
                ;mem[9131] <= 30'b000000001000000000010111010000
                ;mem[9132] <= 30'b000000001000000000010111100000
                ;mem[9133] <= 30'b000000001000000000010111110000
                ;mem[9134] <= 30'b000000001000000000011101010000
                ;mem[9135] <= 30'b000000001000000000011101100000
                ;mem[9136] <= 30'b000000001000000000011101110000
                ;mem[9137] <= 30'b000000001000000000011110000000
                ;mem[9138] <= 30'b000000001000000000011110010000
                ;mem[9139] <= 30'b000000001000000000011110100000
                ;mem[9140] <= 30'b000000001000000000100011110000
                ;mem[9141] <= 30'b000000001000000000100100000000
                ;mem[9142] <= 30'b000000001000000000100100010000
                ;mem[9143] <= 30'b000000001000000000100100100000
                ;mem[9144] <= 30'b000000001000000000100100110000
                ;mem[9145] <= 30'b000000001000000000100101000000
                ;mem[9146] <= 30'b000000001000000000100101010000
                ;mem[9147] <= 30'b000000001000000000100101100000
                ;mem[9148] <= 30'b000000001000000000101010110000
                ;mem[9149] <= 30'b000000001000000000101011000000
                ;mem[9150] <= 30'b000000001000000000101011010000
                ;mem[9151] <= 30'b000000001000000000101011100000
                ;mem[9152] <= 30'b000000001000000000101011110000
                ;mem[9153] <= 30'b000000001000000000101100000000
                ;mem[9154] <= 30'b000000001000000000101100010000
                ;mem[9155] <= 30'b000000001000000000110001010000
                ;mem[9156] <= 30'b000000001000000000110001100000
                ;mem[9157] <= 30'b000000001000000000110001110000
                ;mem[9158] <= 30'b000000001000000000110010000000
                ;mem[9159] <= 30'b000000001000000000110010010000
                ;mem[9160] <= 30'b000000001000000000110010100000
                ;mem[9161] <= 30'b000000001000000000110010110000
                ;mem[9162] <= 30'b000000001000000000110011000000
                ;mem[9163] <= 30'b000000001000000000111000010000
                ;mem[9164] <= 30'b000000001000000000111000100000
                ;mem[9165] <= 30'b000000001000000000111000110000
                ;mem[9166] <= 30'b000000001000000000111001000000
                ;mem[9167] <= 30'b000000001000000000111001010000
                ;mem[9168] <= 30'b000000001000000000111001100000
                ;mem[9169] <= 30'b000000001000000000111001110000
                ;mem[9170] <= 30'b000000001000000000111010000000
                ;mem[9171] <= 30'b000000001000000000111010010000
                ;mem[9172] <= 30'b000000001000000000111111010000
                ;mem[9173] <= 30'b000000001000000000111111100000
                ;mem[9174] <= 30'b000000001000000000111111110000
                ;mem[9175] <= 30'b000000010000000000000000000000
                ;mem[9176] <= 30'b000000010000000000000000010000
                ;mem[9177] <= 30'b000000010000000000000101010000
                ;mem[9178] <= 30'b000000010000000000000101100000
                ;mem[9179] <= 30'b000000010000000000000101110000
                ;mem[9180] <= 30'b000000010000000000000110000000
                ;mem[9181] <= 30'b000000010000000000000110010000
                ;mem[9182] <= 30'b000000010000000000000110100000
                ;mem[9183] <= 30'b000000010000000000000110110000
                ;mem[9184] <= 30'b000000010000000000000111000000
                ;mem[9185] <= 30'b000000010000000000001100010000
                ;mem[9186] <= 30'b000000010000000000001100100000
                ;mem[9187] <= 30'b000000010000000000001100110000
                ;mem[9188] <= 30'b000000010000000000001101000000
                ;mem[9189] <= 30'b000000010000000000001101010000
                ;mem[9190] <= 30'b000000010000000000001101100000
                ;mem[9191] <= 30'b000000010000000000001101110000
                ;mem[9192] <= 30'b000000010000000000001110000000
                ;mem[9193] <= 30'b000000010000000000001110010000
                ;mem[9194] <= 30'b000000010000000000010011010000
                ;mem[9195] <= 30'b000000010000000000010011100000
                ;mem[9196] <= 30'b000000010000000000010011110000
                ;mem[9197] <= 30'b000000010000000000010100000000
                ;mem[9198] <= 30'b000000010000000000010100010000
                ;mem[9199] <= 30'b000000010000000000010100100000
                ;mem[9200] <= 30'b000000010000000000010100110000
                ;mem[9201] <= 30'b000000010000000000010101000000
                ;mem[9202] <= 30'b000000010000000000010101010000
                ;mem[9203] <= 30'b000000010000000000010101100000
                ;mem[9204] <= 30'b000000010000000000011010100000
                ;mem[9205] <= 30'b000000010000000000011010110000
                ;mem[9206] <= 30'b000000010000000000011011000000
                ;mem[9207] <= 30'b000000010000000000011011010000
                ;mem[9208] <= 30'b000000010000000000011011100000
                ;mem[9209] <= 30'b000000010000000000011011110000
                ;mem[9210] <= 30'b000000010000000000011100000000
                ;mem[9211] <= 30'b000000010000000000011100010000
                ;mem[9212] <= 30'b000000010000000000011100100000
                ;mem[9213] <= 30'b000000010000000000011100110000
                ;mem[9214] <= 30'b000000010000000000100011000000
                ;mem[9215] <= 30'b000000010000000000100011010000
                ;mem[9216] <= 30'b000000010000000000100011100000
                ;mem[9217] <= 30'b000000010000000000100011110000
                ;mem[9218] <= 30'b000000010000000000101010000000
                ;mem[9219] <= 30'b000000010000000000101010010000
                ;mem[9220] <= 30'b000000010000000000101010100000
                ;mem[9221] <= 30'b000000010000000000101010110000
                ;mem[9222] <= 30'b000000010000000000110001000000
                ;mem[9223] <= 30'b000000010000000000110001010000
                ;mem[9224] <= 30'b000000010000000000110001100000
                ;mem[9225] <= 30'b000000010000000000110001110000
                ;mem[9226] <= 30'b000000010000000000110110100000
                ;mem[9227] <= 30'b000000010000000000110110110000
                ;mem[9228] <= 30'b000000010000000000110111000000
                ;mem[9229] <= 30'b000000010000000000110111110000
                ;mem[9230] <= 30'b000000010000000000111000000000
                ;mem[9231] <= 30'b000000010000000000111000010000
                ;mem[9232] <= 30'b000000010000000000111000100000
                ;mem[9233] <= 30'b000000010000000000111000110000
                ;mem[9234] <= 30'b000000010000000000111101010000
                ;mem[9235] <= 30'b000000010000000000111101100000
                ;mem[9236] <= 30'b000000010000000000111101110000
                ;mem[9237] <= 30'b000000010000000000111110000000
                ;mem[9238] <= 30'b000000010000000000111110010000
                ;mem[9239] <= 30'b000000010000000000111110100000
                ;mem[9240] <= 30'b000000010000000000111110110000
                ;mem[9241] <= 30'b000000010000000000111111000000
                ;mem[9242] <= 30'b000000010000000000111111010000
                ;mem[9243] <= 30'b000000010000000000111111100000
                ;mem[9244] <= 30'b000000000000000001000101000000
                ;mem[9245] <= 30'b000000000000000001000101010000
                ;mem[9246] <= 30'b000000000000000001000101100000
                ;mem[9247] <= 30'b000000000000000001000101110000
                ;mem[9248] <= 30'b000000000000000001001010100000
                ;mem[9249] <= 30'b000000000000000001001010110000
                ;mem[9250] <= 30'b000000000000000001001011000000
                ;mem[9251] <= 30'b000000000000000001001011110000
                ;mem[9252] <= 30'b000000000000000001001100000000
                ;mem[9253] <= 30'b000000000000000001001100010000
                ;mem[9254] <= 30'b000000000000000001001100100000
                ;mem[9255] <= 30'b000000000000000001001100110000
                ;mem[9256] <= 30'b000000000000000001010001010000
                ;mem[9257] <= 30'b000000000000000001010001100000
                ;mem[9258] <= 30'b000000000000000001010001110000
                ;mem[9259] <= 30'b000000000000000001010010000000
                ;mem[9260] <= 30'b000000000000000001010010010000
                ;mem[9261] <= 30'b000000000000000001010010100000
                ;mem[9262] <= 30'b000000000000000001010010110000
                ;mem[9263] <= 30'b000000000000000001010011000000
                ;mem[9264] <= 30'b000000000000000001010011010000
                ;mem[9265] <= 30'b000000000000000001010011100000
                ;mem[9266] <= 30'b000000000000000001011000100000
                ;mem[9267] <= 30'b000000000000000001011000110000
                ;mem[9268] <= 30'b000000000000000001011001000000
                ;mem[9269] <= 30'b000000000000000001011001010000
                ;mem[9270] <= 30'b000000000000000001011001100000
                ;mem[9271] <= 30'b000000000000000001011001110000
                ;mem[9272] <= 30'b000000000000000001011010000000
                ;mem[9273] <= 30'b000000000000000001011010010000
                ;mem[9274] <= 30'b000000000000000001011010100000
                ;mem[9275] <= 30'b000000000000000001011111100000
                ;mem[9276] <= 30'b000000000000000001011111110000
                ;mem[9277] <= 30'b000000000000000001100000000000
                ;mem[9278] <= 30'b000000000000000001100000010000
                ;mem[9279] <= 30'b000000000000000001100000100000
                ;mem[9280] <= 30'b000000000000000001100000110000
                ;mem[9281] <= 30'b000000000000000001100001000000
                ;mem[9282] <= 30'b000000000000000001100110110000
                ;mem[9283] <= 30'b000000000000000001100111000000
                ;mem[9284] <= 30'b000000000000000001100111010000
                ;mem[9285] <= 30'b000000000000000001100111100000
                ;mem[9286] <= 30'b000000000000000001100111110000
                ;mem[9287] <= 30'b000000000000000000101101000000
                ;mem[9288] <= 30'b000000000000000000101101010000
                ;mem[9289] <= 30'b000000000000000000101101100000
                ;mem[9290] <= 30'b000000000000000000110011100000
                ;mem[9291] <= 30'b000000000000000000110011110000
                ;mem[9292] <= 30'b000000000000000000110100000000
                ;mem[9293] <= 30'b000000000000000000110100010000
                ;mem[9294] <= 30'b000000000000000000110100100000
                ;mem[9295] <= 30'b000000000000000000110100110000
                ;mem[9296] <= 30'b000000000000000000110101000000
                ;mem[9297] <= 30'b000000000000000000110101010000
                ;mem[9298] <= 30'b000000000000000000110101100000
                ;mem[9299] <= 30'b000000000000000000110101110000
                ;mem[9300] <= 30'b000000000000000000110110000000
                ;mem[9301] <= 30'b000000000000000000110110010000
                ;mem[9302] <= 30'b000000000000000000111010010000
                ;mem[9303] <= 30'b000000000000000000111010100000
                ;mem[9304] <= 30'b000000000000000000111010110000
                ;mem[9305] <= 30'b000000000000000000111011000000
                ;mem[9306] <= 30'b000000000000000000111011010000
                ;mem[9307] <= 30'b000000000000000000111011100000
                ;mem[9308] <= 30'b000000000000000000111011110000
                ;mem[9309] <= 30'b000000000000000000111100000000
                ;mem[9310] <= 30'b000000000000000000111100010000
                ;mem[9311] <= 30'b000000000000000000111100100000
                ;mem[9312] <= 30'b000000000000000000111100110000
                ;mem[9313] <= 30'b000000000000000000111101000000
                ;mem[9314] <= 30'b000000000000000000111101010000
                ;mem[9315] <= 30'b000000000000000000111101100000
                ;mem[9316] <= 30'b000000001000000000000001000000
                ;mem[9317] <= 30'b000000001000000000000001010000
                ;mem[9318] <= 30'b000000001000000000000001100000
                ;mem[9319] <= 30'b000000001000000000000111100000
                ;mem[9320] <= 30'b000000001000000000000111110000
                ;mem[9321] <= 30'b000000001000000000001000000000
                ;mem[9322] <= 30'b000000001000000000001000010000
                ;mem[9323] <= 30'b000000001000000000001000100000
                ;mem[9324] <= 30'b000000001000000000001000110000
                ;mem[9325] <= 30'b000000001000000000001001000000
                ;mem[9326] <= 30'b000000001000000000001001010000
                ;mem[9327] <= 30'b000000001000000000001001100000
                ;mem[9328] <= 30'b000000001000000000001001110000
                ;mem[9329] <= 30'b000000001000000000001010000000
                ;mem[9330] <= 30'b000000001000000000001010010000
                ;mem[9331] <= 30'b000000001000000000001110010000
                ;mem[9332] <= 30'b000000001000000000001110100000
                ;mem[9333] <= 30'b000000001000000000001110110000
                ;mem[9334] <= 30'b000000001000000000001111000000
                ;mem[9335] <= 30'b000000001000000000001111010000
                ;mem[9336] <= 30'b000000001000000000001111100000
                ;mem[9337] <= 30'b000000001000000000001111110000
                ;mem[9338] <= 30'b000000001000000000010000000000
                ;mem[9339] <= 30'b000000001000000000010000010000
                ;mem[9340] <= 30'b000000001000000000010000100000
                ;mem[9341] <= 30'b000000001000000000010000110000
                ;mem[9342] <= 30'b000000001000000000010001000000
                ;mem[9343] <= 30'b000000001000000000010001010000
                ;mem[9344] <= 30'b000000001000000000010001100000
                ;mem[9345] <= 30'b000000001000000000010101000000
                ;mem[9346] <= 30'b000000001000000000010101010000
                ;mem[9347] <= 30'b000000001000000000010101100000
                ;mem[9348] <= 30'b000000001000000000010101110000
                ;mem[9349] <= 30'b000000001000000000010110010000
                ;mem[9350] <= 30'b000000001000000000010110100000
                ;mem[9351] <= 30'b000000001000000000011000010000
                ;mem[9352] <= 30'b000000001000000000011000100000
                ;mem[9353] <= 30'b000000001000000000011000110000
                ;mem[9354] <= 30'b000000001000000000011011110000
                ;mem[9355] <= 30'b000000001000000000011100000000
                ;mem[9356] <= 30'b000000001000000000011100010000
                ;mem[9357] <= 30'b000000001000000000011111100000
                ;mem[9358] <= 30'b000000001000000000011111110000
                ;mem[9359] <= 30'b000000001000000000100010110000
                ;mem[9360] <= 30'b000000001000000000100011000000
                ;mem[9361] <= 30'b000000001000000000100110110000
                ;mem[9362] <= 30'b000000001000000000100111000000
                ;mem[9363] <= 30'b000000001000000000101001100000
                ;mem[9364] <= 30'b000000001000000000101001110000
                ;mem[9365] <= 30'b000000001000000000101101110000
                ;mem[9366] <= 30'b000000001000000000101110000000
                ;mem[9367] <= 30'b000000001000000000110000010000
                ;mem[9368] <= 30'b000000001000000000110000100000
                ;mem[9369] <= 30'b000000001000000000110000110000
                ;mem[9370] <= 30'b000000001000000000110100110000
                ;mem[9371] <= 30'b000000001000000000110101000000
                ;mem[9372] <= 30'b000000001000000000110111010000
                ;mem[9373] <= 30'b000000001000000000110111100000
                ;mem[9374] <= 30'b000000001000000000111011110000
                ;mem[9375] <= 30'b000000001000000000111100000000
                ;mem[9376] <= 30'b000000001000000000111110010000
                ;mem[9377] <= 30'b000000001000000000111110100000
                ;mem[9378] <= 30'b000000010000000000000001110000
                ;mem[9379] <= 30'b000000010000000000000010000000
                ;mem[9380] <= 30'b000000010000000000000100010000
                ;mem[9381] <= 30'b000000010000000000000100100000
                ;mem[9382] <= 30'b000000010000000000000100110000
                ;mem[9383] <= 30'b000000010000000000001000110000
                ;mem[9384] <= 30'b000000010000000000001001000000
                ;mem[9385] <= 30'b000000010000000000001011010000
                ;mem[9386] <= 30'b000000010000000000001011100000
                ;mem[9387] <= 30'b000000010000000000001111110000
                ;mem[9388] <= 30'b000000010000000000010000000000
                ;mem[9389] <= 30'b000000010000000000010010010000
                ;mem[9390] <= 30'b000000010000000000010010100000
                ;mem[9391] <= 30'b000000010000000000010110100000
                ;mem[9392] <= 30'b000000010000000000010110110000
                ;mem[9393] <= 30'b000000010000000000010111000000
                ;mem[9394] <= 30'b000000010000000000011001010000
                ;mem[9395] <= 30'b000000010000000000011001100000
                ;mem[9396] <= 30'b000000010000000000011101100000
                ;mem[9397] <= 30'b000000010000000000011101110000
                ;mem[9398] <= 30'b000000010000000000011110000000
                ;mem[9399] <= 30'b000000010000000000100000010000
                ;mem[9400] <= 30'b000000010000000000100000100000
                ;mem[9401] <= 30'b000000010000000000100100010000
                ;mem[9402] <= 30'b000000010000000000100100100000
                ;mem[9403] <= 30'b000000010000000000100100110000
                ;mem[9404] <= 30'b000000010000000000100111010000
                ;mem[9405] <= 30'b000000010000000000100111100000
                ;mem[9406] <= 30'b000000010000000000100111110000
                ;mem[9407] <= 30'b000000010000000000101010110000
                ;mem[9408] <= 30'b000000010000000000101011000000
                ;mem[9409] <= 30'b000000010000000000101011010000
                ;mem[9410] <= 30'b000000010000000000101011100000
                ;mem[9411] <= 30'b000000010000000000101110100000
                ;mem[9412] <= 30'b000000010000000000101110110000
                ;mem[9413] <= 30'b000000010000000000101111000000
                ;mem[9414] <= 30'b000000010000000000101111010000
                ;mem[9415] <= 30'b000000010000000000101111100000
                ;mem[9416] <= 30'b000000010000000000110000010000
                ;mem[9417] <= 30'b000000010000000000110000100000
                ;mem[9418] <= 30'b000000010000000000110000110000
                ;mem[9419] <= 30'b000000010000000000110001000000
                ;mem[9420] <= 30'b000000010000000000110001010000
                ;mem[9421] <= 30'b000000010000000000110001100000
                ;mem[9422] <= 30'b000000010000000000110001110000
                ;mem[9423] <= 30'b000000010000000000110010000000
                ;mem[9424] <= 30'b000000010000000000110010010000
                ;mem[9425] <= 30'b000000010000000000110101110000
                ;mem[9426] <= 30'b000000010000000000110110000000
                ;mem[9427] <= 30'b000000010000000000110110010000
                ;mem[9428] <= 30'b000000010000000000110110100000
                ;mem[9429] <= 30'b000000010000000000110110110000
                ;mem[9430] <= 30'b000000010000000000110111000000
                ;mem[9431] <= 30'b000000010000000000110111010000
                ;mem[9432] <= 30'b000000010000000000110111100000
                ;mem[9433] <= 30'b000000010000000000110111110000
                ;mem[9434] <= 30'b000000010000000000111000000000
                ;mem[9435] <= 30'b000000010000000000111000010000
                ;mem[9436] <= 30'b000000010000000000111000100000
                ;mem[9437] <= 30'b000000010000000000111101010000
                ;mem[9438] <= 30'b000000010000000000111101100000
                ;mem[9439] <= 30'b000000010000000000111101110000
                ;mem[9440] <= 30'b000000010000000000111110000000
                ;mem[9441] <= 30'b000000010000000000111110010000
                ;mem[9442] <= 30'b000000010000000000111110100000
                ;mem[9443] <= 30'b000000010000000000111110110000
                ;mem[9444] <= 30'b000000000000000001000010100000
                ;mem[9445] <= 30'b000000000000000001000010110000
                ;mem[9446] <= 30'b000000000000000001000011000000
                ;mem[9447] <= 30'b000000000000000001000011010000
                ;mem[9448] <= 30'b000000000000000001000011100000
                ;mem[9449] <= 30'b000000000000000001000100010000
                ;mem[9450] <= 30'b000000000000000001000100100000
                ;mem[9451] <= 30'b000000000000000001000100110000
                ;mem[9452] <= 30'b000000000000000001000101000000
                ;mem[9453] <= 30'b000000000000000001000101010000
                ;mem[9454] <= 30'b000000000000000001000101100000
                ;mem[9455] <= 30'b000000000000000001000101110000
                ;mem[9456] <= 30'b000000000000000001000110000000
                ;mem[9457] <= 30'b000000000000000001000110010000
                ;mem[9458] <= 30'b000000000000000001001001110000
                ;mem[9459] <= 30'b000000000000000001001010000000
                ;mem[9460] <= 30'b000000000000000001001010010000
                ;mem[9461] <= 30'b000000000000000001001010100000
                ;mem[9462] <= 30'b000000000000000001001010110000
                ;mem[9463] <= 30'b000000000000000001001011000000
                ;mem[9464] <= 30'b000000000000000001001011010000
                ;mem[9465] <= 30'b000000000000000001001011100000
                ;mem[9466] <= 30'b000000000000000001001011110000
                ;mem[9467] <= 30'b000000000000000001001100000000
                ;mem[9468] <= 30'b000000000000000001001100010000
                ;mem[9469] <= 30'b000000000000000001001100100000
                ;mem[9470] <= 30'b000000000000000001010001010000
                ;mem[9471] <= 30'b000000000000000001010001100000
                ;mem[9472] <= 30'b000000000000000001010001110000
                ;mem[9473] <= 30'b000000000000000001010010000000
                ;mem[9474] <= 30'b000000000000000001010010010000
                ;mem[9475] <= 30'b000000000000000001010010100000
                ;mem[9476] <= 30'b000000000000000001010010110000
                ;mem[9477] <= 30'b000000000000000000111000100000
                ;mem[9478] <= 30'b000000000000000000111000110000
                ;mem[9479] <= 30'b000000000000000000111001000000
                ;mem[9480] <= 30'b000000000000000000111001010000
                ;mem[9481] <= 30'b000000000000000000111001100000
                ;mem[9482] <= 30'b000000000000000000111001110000
                ;mem[9483] <= 30'b000000000000000000111010000000
                ;mem[9484] <= 30'b000000000000000000111010010000
                ;mem[9485] <= 30'b000000000000000000111010100000
                ;mem[9486] <= 30'b000000000000000000111010110000
                ;mem[9487] <= 30'b000000000000000000111011000000
                ;mem[9488] <= 30'b000000000000000000111011010000
                ;mem[9489] <= 30'b000000000000000000111011100000
                ;mem[9490] <= 30'b000000000000000000111011110000
                ;mem[9491] <= 30'b000000000000000000111100000000
                ;mem[9492] <= 30'b000000000000000000111111100000
                ;mem[9493] <= 30'b000000000000000000111111110000
                ;mem[9494] <= 30'b000000001000000000001100100000
                ;mem[9495] <= 30'b000000001000000000001100110000
                ;mem[9496] <= 30'b000000001000000000001101000000
                ;mem[9497] <= 30'b000000001000000000001101010000
                ;mem[9498] <= 30'b000000001000000000001101100000
                ;mem[9499] <= 30'b000000001000000000001101110000
                ;mem[9500] <= 30'b000000001000000000001110000000
                ;mem[9501] <= 30'b000000001000000000001110010000
                ;mem[9502] <= 30'b000000001000000000001110100000
                ;mem[9503] <= 30'b000000001000000000001110110000
                ;mem[9504] <= 30'b000000001000000000001111000000
                ;mem[9505] <= 30'b000000001000000000001111010000
                ;mem[9506] <= 30'b000000001000000000001111100000
                ;mem[9507] <= 30'b000000001000000000001111110000
                ;mem[9508] <= 30'b000000001000000000010000000000
                ;mem[9509] <= 30'b000000001000000000010011100000
                ;mem[9510] <= 30'b000000001000000000010011110000
                ;mem[9511] <= 30'b000000001000000000010100000000
                ;mem[9512] <= 30'b000000001000000000010100010000
                ;mem[9513] <= 30'b000000001000000000010100100000
                ;mem[9514] <= 30'b000000001000000000010100110000
                ;mem[9515] <= 30'b000000001000000000010101000000
                ;mem[9516] <= 30'b000000001000000000010101010000
                ;mem[9517] <= 30'b000000001000000000010101100000
                ;mem[9518] <= 30'b000000001000000000010101110000
                ;mem[9519] <= 30'b000000001000000000010110000000
                ;mem[9520] <= 30'b000000001000000000010110010000
                ;mem[9521] <= 30'b000000001000000000010110100000
                ;mem[9522] <= 30'b000000001000000000010110110000
                ;mem[9523] <= 30'b000000001000000000010111000000
                ;mem[9524] <= 30'b000000001000000000010111010000
                ;mem[9525] <= 30'b000000001000000000010111100000
                ;mem[9526] <= 30'b000000001000000000010111110000
                ;mem[9527] <= 30'b000000001000000000011101000000
                ;mem[9528] <= 30'b000000001000000000011101100000
                ;mem[9529] <= 30'b000000001000000000011101110000
                ;mem[9530] <= 30'b000000001000000000011110000000
                ;mem[9531] <= 30'b000000001000000000011110010000
                ;mem[9532] <= 30'b000000001000000000011110100000
                ;mem[9533] <= 30'b000000001000000000011110110000
                ;mem[9534] <= 30'b000000001000000000011111000000
                ;mem[9535] <= 30'b000000001000000000100101010000
                ;mem[9536] <= 30'b000000001000000000100101100000
                ;mem[9537] <= 30'b000000001000000000100101110000
                ;mem[9538] <= 30'b000000001000000000100110000000
                ;mem[9539] <= 30'b000000001000000000100110010000
                ;mem[9540] <= 30'b000000001000000000101100110000
                ;mem[9541] <= 30'b000000001000000000101101000000
                ;mem[9542] <= 30'b000000001000000000101101010000
                ;mem[9543] <= 30'b000000001000000000110011110000
                ;mem[9544] <= 30'b000000001000000000110100000000
                ;mem[9545] <= 30'b000000001000000000110100010000
                ;mem[9546] <= 30'b000000001000000000111010100000
                ;mem[9547] <= 30'b000000001000000000111010110000
                ;mem[9548] <= 30'b000000001000000000111011000000
                ;mem[9549] <= 30'b000000010000000000000000110000
                ;mem[9550] <= 30'b000000010000000000000001000000
                ;mem[9551] <= 30'b000000010000000000000001010000
                ;mem[9552] <= 30'b000000010000000000000111110000
                ;mem[9553] <= 30'b000000010000000000001000000000
                ;mem[9554] <= 30'b000000010000000000001000010000
                ;mem[9555] <= 30'b000000010000000000001110100000
                ;mem[9556] <= 30'b000000010000000000001110110000
                ;mem[9557] <= 30'b000000010000000000001111000000
                ;mem[9558] <= 30'b000000010000000000010101100000
                ;mem[9559] <= 30'b000000010000000000010101110000
                ;mem[9560] <= 30'b000000010000000000010110000000
                ;mem[9561] <= 30'b000000010000000000011100010000
                ;mem[9562] <= 30'b000000010000000000011100100000
                ;mem[9563] <= 30'b000000010000000000011100110000
                ;mem[9564] <= 30'b000000010000000000100011000000
                ;mem[9565] <= 30'b000000010000000000100011010000
                ;mem[9566] <= 30'b000000010000000000100011100000
                ;mem[9567] <= 30'b000000010000000000101001110000
                ;mem[9568] <= 30'b000000010000000000101010000000
                ;mem[9569] <= 30'b000000010000000000101010010000
                ;mem[9570] <= 30'b000000010000000000110000100000
                ;mem[9571] <= 30'b000000010000000000110000110000
                ;mem[9572] <= 30'b000000010000000000110001000000
                ;mem[9573] <= 30'b000000010000000000110001010000
                ;mem[9574] <= 30'b000000010000000000110111100000
                ;mem[9575] <= 30'b000000010000000000110111110000
                ;mem[9576] <= 30'b000000010000000000111000000000
                ;mem[9577] <= 30'b000000010000000000111110010000
                ;mem[9578] <= 30'b000000010000000000111110100000
                ;mem[9579] <= 30'b000000010000000000111110110000
                ;mem[9580] <= 30'b000000000000000001000100100000
                ;mem[9581] <= 30'b000000000000000001000100110000
                ;mem[9582] <= 30'b000000000000000001000101000000
                ;mem[9583] <= 30'b000000000000000001000101010000
                ;mem[9584] <= 30'b000000000000000001001011100000
                ;mem[9585] <= 30'b000000000000000001001011110000
                ;mem[9586] <= 30'b000000000000000001001100000000
                ;mem[9587] <= 30'b000000000000000001010010010000
                ;mem[9588] <= 30'b000000000000000001010010100000
                ;mem[9589] <= 30'b000000000000000001010010110000
                ;mem[9590] <= 30'b000000000000000001011001000000
                ;mem[9591] <= 30'b000000000000000001011001010000
                ;mem[9592] <= 30'b000000000000000001011001100000
                ;mem[9593] <= 30'b000000000000000001011111110000
                ;mem[9594] <= 30'b000000000000000001100000000000
                ;mem[9595] <= 30'b000000000000000001100000010000
                ;mem[9596] <= 30'b000000000000000001100000100000
                ;mem[9597] <= 30'b000000000000000001100110110000
                ;mem[9598] <= 30'b000000000000000001100111000000
                ;mem[9599] <= 30'b000000000000000001100111010000
                ;mem[9600] <= 30'b000000000000000001101101100000
                ;mem[9601] <= 30'b000000000000000001101101110000
                ;mem[9602] <= 30'b000000000000000001101110000000
                ;mem[9603] <= 30'b000000000000000000011111000000
                ;mem[9604] <= 30'b000000000000000000011111010000
                ;mem[9605] <= 30'b000000000000000000011111100000
                ;mem[9606] <= 30'b000000000000000000011111110000
                ;mem[9607] <= 30'b000000000000000000100000000000
                ;mem[9608] <= 30'b000000000000000000100101110000
                ;mem[9609] <= 30'b000000000000000000100110000000
                ;mem[9610] <= 30'b000000000000000000100110010000
                ;mem[9611] <= 30'b000000000000000000100110100000
                ;mem[9612] <= 30'b000000000000000000100110110000
                ;mem[9613] <= 30'b000000000000000000100111000000
                ;mem[9614] <= 30'b000000000000000000100111010000
                ;mem[9615] <= 30'b000000000000000000100111100000
                ;mem[9616] <= 30'b000000000000000000101100100000
                ;mem[9617] <= 30'b000000000000000000101100110000
                ;mem[9618] <= 30'b000000000000000000101101000000
                ;mem[9619] <= 30'b000000000000000000101101010000
                ;mem[9620] <= 30'b000000000000000000101101100000
                ;mem[9621] <= 30'b000000000000000000101101110000
                ;mem[9622] <= 30'b000000000000000000101110000000
                ;mem[9623] <= 30'b000000000000000000101110010000
                ;mem[9624] <= 30'b000000000000000000101110100000
                ;mem[9625] <= 30'b000000000000000000101110110000
                ;mem[9626] <= 30'b000000000000000000101111000000
                ;mem[9627] <= 30'b000000000000000000110011010000
                ;mem[9628] <= 30'b000000000000000000110011100000
                ;mem[9629] <= 30'b000000000000000000110011110000
                ;mem[9630] <= 30'b000000000000000000110100000000
                ;mem[9631] <= 30'b000000000000000000110100010000
                ;mem[9632] <= 30'b000000000000000000110101000000
                ;mem[9633] <= 30'b000000000000000000110101010000
                ;mem[9634] <= 30'b000000000000000000110101100000
                ;mem[9635] <= 30'b000000000000000000110101110000
                ;mem[9636] <= 30'b000000000000000000110110000000
                ;mem[9637] <= 30'b000000000000000000110110010000
                ;mem[9638] <= 30'b000000000000000000111010010000
                ;mem[9639] <= 30'b000000000000000000111010100000
                ;mem[9640] <= 30'b000000000000000000111010110000
                ;mem[9641] <= 30'b000000000000000000111011000000
                ;mem[9642] <= 30'b000000000000000000111100100000
                ;mem[9643] <= 30'b000000000000000000111100110000
                ;mem[9644] <= 30'b000000000000000000111101000000
                ;mem[9645] <= 30'b000000000000000000111101010000
                ;mem[9646] <= 30'b000000000000000000111101100000
                ;mem[9647] <= 30'b000000001000000000000000100000
                ;mem[9648] <= 30'b000000001000000000000000110000
                ;mem[9649] <= 30'b000000001000000000000001000000
                ;mem[9650] <= 30'b000000001000000000000001010000
                ;mem[9651] <= 30'b000000001000000000000001100000
                ;mem[9652] <= 30'b000000001000000000000001110000
                ;mem[9653] <= 30'b000000001000000000000010000000
                ;mem[9654] <= 30'b000000001000000000000010010000
                ;mem[9655] <= 30'b000000001000000000000010100000
                ;mem[9656] <= 30'b000000001000000000000010110000
                ;mem[9657] <= 30'b000000001000000000000011000000
                ;mem[9658] <= 30'b000000001000000000000111010000
                ;mem[9659] <= 30'b000000001000000000000111100000
                ;mem[9660] <= 30'b000000001000000000000111110000
                ;mem[9661] <= 30'b000000001000000000001000000000
                ;mem[9662] <= 30'b000000001000000000001000010000
                ;mem[9663] <= 30'b000000001000000000001001000000
                ;mem[9664] <= 30'b000000001000000000001001010000
                ;mem[9665] <= 30'b000000001000000000001001100000
                ;mem[9666] <= 30'b000000001000000000001001110000
                ;mem[9667] <= 30'b000000001000000000001010000000
                ;mem[9668] <= 30'b000000001000000000001010010000
                ;mem[9669] <= 30'b000000001000000000001110010000
                ;mem[9670] <= 30'b000000001000000000001110100000
                ;mem[9671] <= 30'b000000001000000000001110110000
                ;mem[9672] <= 30'b000000001000000000001111000000
                ;mem[9673] <= 30'b000000001000000000010000100000
                ;mem[9674] <= 30'b000000001000000000010000110000
                ;mem[9675] <= 30'b000000001000000000010001000000
                ;mem[9676] <= 30'b000000001000000000010001010000
                ;mem[9677] <= 30'b000000001000000000010001100000
                ;mem[9678] <= 30'b000000001000000000010101000000
                ;mem[9679] <= 30'b000000001000000000010101010000
                ;mem[9680] <= 30'b000000001000000000010101100000
                ;mem[9681] <= 30'b000000001000000000010101110000
                ;mem[9682] <= 30'b000000001000000000010111110000
                ;mem[9683] <= 30'b000000001000000000011000000000
                ;mem[9684] <= 30'b000000001000000000011000010000
                ;mem[9685] <= 30'b000000001000000000011000100000
                ;mem[9686] <= 30'b000000001000000000011011110000
                ;mem[9687] <= 30'b000000001000000000011100000000
                ;mem[9688] <= 30'b000000001000000000011100010000
                ;mem[9689] <= 30'b000000001000000000011100100000
                ;mem[9690] <= 30'b000000001000000000011100110000
                ;mem[9691] <= 30'b000000001000000000011111000000
                ;mem[9692] <= 30'b000000001000000000011111010000
                ;mem[9693] <= 30'b000000001000000000011111100000
                ;mem[9694] <= 30'b000000001000000000100010110000
                ;mem[9695] <= 30'b000000001000000000100011000000
                ;mem[9696] <= 30'b000000001000000000100011010000
                ;mem[9697] <= 30'b000000001000000000100011100000
                ;mem[9698] <= 30'b000000001000000000100110000000
                ;mem[9699] <= 30'b000000001000000000100110010000
                ;mem[9700] <= 30'b000000001000000000100110100000
                ;mem[9701] <= 30'b000000001000000000101001110000
                ;mem[9702] <= 30'b000000001000000000101010000000
                ;mem[9703] <= 30'b000000001000000000101010010000
                ;mem[9704] <= 30'b000000001000000000101101000000
                ;mem[9705] <= 30'b000000001000000000101101010000
                ;mem[9706] <= 30'b000000001000000000101101100000
                ;mem[9707] <= 30'b000000001000000000110000100000
                ;mem[9708] <= 30'b000000001000000000110000110000
                ;mem[9709] <= 30'b000000001000000000110001000000
                ;mem[9710] <= 30'b000000001000000000110001010000
                ;mem[9711] <= 30'b000000001000000000110100000000
                ;mem[9712] <= 30'b000000001000000000110100010000
                ;mem[9713] <= 30'b000000001000000000110100100000
                ;mem[9714] <= 30'b000000001000000000110100110000
                ;mem[9715] <= 30'b000000001000000000110111100000
                ;mem[9716] <= 30'b000000001000000000110111110000
                ;mem[9717] <= 30'b000000001000000000111000000000
                ;mem[9718] <= 30'b000000001000000000111011000000
                ;mem[9719] <= 30'b000000001000000000111011010000
                ;mem[9720] <= 30'b000000001000000000111011100000
                ;mem[9721] <= 30'b000000001000000000111011110000
                ;mem[9722] <= 30'b000000001000000000111110100000
                ;mem[9723] <= 30'b000000001000000000111110110000
                ;mem[9724] <= 30'b000000001000000000111111000000
                ;mem[9725] <= 30'b000000010000000000000001000000
                ;mem[9726] <= 30'b000000010000000000000001010000
                ;mem[9727] <= 30'b000000010000000000000001100000
                ;mem[9728] <= 30'b000000010000000000000100100000
                ;mem[9729] <= 30'b000000010000000000000100110000
                ;mem[9730] <= 30'b000000010000000000000101000000
                ;mem[9731] <= 30'b000000010000000000000101010000
                ;mem[9732] <= 30'b000000010000000000001000000000
                ;mem[9733] <= 30'b000000010000000000001000010000
                ;mem[9734] <= 30'b000000010000000000001000100000
                ;mem[9735] <= 30'b000000010000000000001000110000
                ;mem[9736] <= 30'b000000010000000000001011100000
                ;mem[9737] <= 30'b000000010000000000001011110000
                ;mem[9738] <= 30'b000000010000000000001100000000
                ;mem[9739] <= 30'b000000010000000000001111000000
                ;mem[9740] <= 30'b000000010000000000001111010000
                ;mem[9741] <= 30'b000000010000000000001111100000
                ;mem[9742] <= 30'b000000010000000000001111110000
                ;mem[9743] <= 30'b000000010000000000010010100000
                ;mem[9744] <= 30'b000000010000000000010010110000
                ;mem[9745] <= 30'b000000010000000000010011000000
                ;mem[9746] <= 30'b000000010000000000010110000000
                ;mem[9747] <= 30'b000000010000000000010110010000
                ;mem[9748] <= 30'b000000010000000000010110100000
                ;mem[9749] <= 30'b000000010000000000010110110000
                ;mem[9750] <= 30'b000000010000000000011001100000
                ;mem[9751] <= 30'b000000010000000000011001110000
                ;mem[9752] <= 30'b000000010000000000011010000000
                ;mem[9753] <= 30'b000000010000000000011010010000
                ;mem[9754] <= 30'b000000010000000000011101000000
                ;mem[9755] <= 30'b000000010000000000011101010000
                ;mem[9756] <= 30'b000000010000000000011101100000
                ;mem[9757] <= 30'b000000010000000000100000100000
                ;mem[9758] <= 30'b000000010000000000100000110000
                ;mem[9759] <= 30'b000000010000000000100001000000
                ;mem[9760] <= 30'b000000010000000000100001010000
                ;mem[9761] <= 30'b000000010000000000100011110000
                ;mem[9762] <= 30'b000000010000000000100100000000
                ;mem[9763] <= 30'b000000010000000000100100010000
                ;mem[9764] <= 30'b000000010000000000100100100000
                ;mem[9765] <= 30'b000000010000000000100111110000
                ;mem[9766] <= 30'b000000010000000000101000000000
                ;mem[9767] <= 30'b000000010000000000101000010000
                ;mem[9768] <= 30'b000000010000000000101010110000
                ;mem[9769] <= 30'b000000010000000000101011000000
                ;mem[9770] <= 30'b000000010000000000101011010000
                ;mem[9771] <= 30'b000000010000000000101011100000
                ;mem[9772] <= 30'b000000010000000000101110110000
                ;mem[9773] <= 30'b000000010000000000101111000000
                ;mem[9774] <= 30'b000000010000000000101111010000
                ;mem[9775] <= 30'b000000010000000000110001010000
                ;mem[9776] <= 30'b000000010000000000110001100000
                ;mem[9777] <= 30'b000000010000000000110001110000
                ;mem[9778] <= 30'b000000010000000000110010000000
                ;mem[9779] <= 30'b000000010000000000110010010000
                ;mem[9780] <= 30'b000000010000000000110010100000
                ;mem[9781] <= 30'b000000010000000000110101110000
                ;mem[9782] <= 30'b000000010000000000110110000000
                ;mem[9783] <= 30'b000000010000000000110110010000
                ;mem[9784] <= 30'b000000010000000000110110100000
                ;mem[9785] <= 30'b000000010000000000110111000000
                ;mem[9786] <= 30'b000000010000000000110111010000
                ;mem[9787] <= 30'b000000010000000000110111100000
                ;mem[9788] <= 30'b000000010000000000110111110000
                ;mem[9789] <= 30'b000000010000000000111000000000
                ;mem[9790] <= 30'b000000010000000000111000010000
                ;mem[9791] <= 30'b000000010000000000111000100000
                ;mem[9792] <= 30'b000000010000000000111000110000
                ;mem[9793] <= 30'b000000010000000000111001000000
                ;mem[9794] <= 30'b000000010000000000111001010000
                ;mem[9795] <= 30'b000000010000000000111101000000
                ;mem[9796] <= 30'b000000010000000000111101010000
                ;mem[9797] <= 30'b000000010000000000111101100000
                ;mem[9798] <= 30'b000000010000000000111101110000
                ;mem[9799] <= 30'b000000010000000000111110000000
                ;mem[9800] <= 30'b000000010000000000111110010000
                ;mem[9801] <= 30'b000000010000000000111110100000
                ;mem[9802] <= 30'b000000010000000000111110110000
                ;mem[9803] <= 30'b000000010000000000111111000000
                ;mem[9804] <= 30'b000000010000000000111111010000
                ;mem[9805] <= 30'b000000010000000000111111100000
                ;mem[9806] <= 30'b000000010000000000111111110000
                ;mem[9807] <= 30'b000000000000000001000010110000
                ;mem[9808] <= 30'b000000000000000001000011000000
                ;mem[9809] <= 30'b000000000000000001000011010000
                ;mem[9810] <= 30'b000000000000000001000101010000
                ;mem[9811] <= 30'b000000000000000001000101100000
                ;mem[9812] <= 30'b000000000000000001000101110000
                ;mem[9813] <= 30'b000000000000000001000110000000
                ;mem[9814] <= 30'b000000000000000001000110010000
                ;mem[9815] <= 30'b000000000000000001000110100000
                ;mem[9816] <= 30'b000000000000000001001001110000
                ;mem[9817] <= 30'b000000000000000001001010000000
                ;mem[9818] <= 30'b000000000000000001001010010000
                ;mem[9819] <= 30'b000000000000000001001010100000
                ;mem[9820] <= 30'b000000000000000001001011000000
                ;mem[9821] <= 30'b000000000000000001001011010000
                ;mem[9822] <= 30'b000000000000000001001011100000
                ;mem[9823] <= 30'b000000000000000001001011110000
                ;mem[9824] <= 30'b000000000000000001001100000000
                ;mem[9825] <= 30'b000000000000000001001100010000
                ;mem[9826] <= 30'b000000000000000001001100100000
                ;mem[9827] <= 30'b000000000000000001001100110000
                ;mem[9828] <= 30'b000000000000000001001101000000
                ;mem[9829] <= 30'b000000000000000001001101010000
                ;mem[9830] <= 30'b000000000000000001010001000000
                ;mem[9831] <= 30'b000000000000000001010001010000
                ;mem[9832] <= 30'b000000000000000001010001100000
                ;mem[9833] <= 30'b000000000000000001010001110000
                ;mem[9834] <= 30'b000000000000000001010010000000
                ;mem[9835] <= 30'b000000000000000001010010010000
                ;mem[9836] <= 30'b000000000000000001010010100000
                ;mem[9837] <= 30'b000000000000000001010010110000
                ;mem[9838] <= 30'b000000000000000001010011000000
                ;mem[9839] <= 30'b000000000000000001010011010000
                ;mem[9840] <= 30'b000000000000000001010011100000
                ;mem[9841] <= 30'b000000000000000001010011110000
                ;mem[9842] <= 30'b000000000000000001010100000000
                ;mem[9843] <= 30'b000000000000000001011000000000
                ;mem[9844] <= 30'b000000000000000001011000010000
                ;mem[9845] <= 30'b000000000000000001011000100000
                ;mem[9846] <= 30'b000000000000000001011000110000
                ;mem[9847] <= 30'b000000000000000001011001000000
                ;mem[9848] <= 30'b000000000000000001011001010000
                ;mem[9849] <= 30'b000000000000000001011001100000
                ;mem[9850] <= 30'b000000000000000001011001110000
                ;mem[9851] <= 30'b000000000000000001011010000000
                ;mem[9852] <= 30'b000000000000000001011010010000
                ;mem[9853] <= 30'b000000000000000001011010100000
                ;mem[9854] <= 30'b000000000000000001011111010000
                ;mem[9855] <= 30'b000000000000000001011111100000
                ;mem[9856] <= 30'b000000000000000001011111110000
                ;mem[9857] <= 30'b000000000000000000011110000000
                ;mem[9858] <= 30'b000000000000000000011110010000
                ;mem[9859] <= 30'b000000000000000000011110100000
                ;mem[9860] <= 30'b000000000000000000011110110000
                ;mem[9861] <= 30'b000000000000000000011111000000
                ;mem[9862] <= 30'b000000000000000000011111010000
                ;mem[9863] <= 30'b000000000000000000011111100000
                ;mem[9864] <= 30'b000000000000000000011111110000
                ;mem[9865] <= 30'b000000000000000000100000000000
                ;mem[9866] <= 30'b000000000000000000100000010000
                ;mem[9867] <= 30'b000000000000000000100100110000
                ;mem[9868] <= 30'b000000000000000000100101000000
                ;mem[9869] <= 30'b000000000000000000100101010000
                ;mem[9870] <= 30'b000000000000000000100101100000
                ;mem[9871] <= 30'b000000000000000000100101110000
                ;mem[9872] <= 30'b000000000000000000100110000000
                ;mem[9873] <= 30'b000000000000000000100110010000
                ;mem[9874] <= 30'b000000000000000000100110100000
                ;mem[9875] <= 30'b000000000000000000100110110000
                ;mem[9876] <= 30'b000000000000000000100111000000
                ;mem[9877] <= 30'b000000000000000000100111010000
                ;mem[9878] <= 30'b000000000000000000100111100000
                ;mem[9879] <= 30'b000000000000000000101011110000
                ;mem[9880] <= 30'b000000000000000000101100000000
                ;mem[9881] <= 30'b000000000000000000101100010000
                ;mem[9882] <= 30'b000000000000000000101100100000
                ;mem[9883] <= 30'b000000000000000000101100110000
                ;mem[9884] <= 30'b000000000000000000101110010000
                ;mem[9885] <= 30'b000000000000000000101110100000
                ;mem[9886] <= 30'b000000000000000000101110110000
                ;mem[9887] <= 30'b000000000000000000110011000000
                ;mem[9888] <= 30'b000000000000000000110011010000
                ;mem[9889] <= 30'b000000000000000000110101100000
                ;mem[9890] <= 30'b000000000000000000110101110000
                ;mem[9891] <= 30'b000000000000000000110110000000
                ;mem[9892] <= 30'b000000000000000000111100110000
                ;mem[9893] <= 30'b000000000000000000111101000000
                ;mem[9894] <= 30'b000000001000000000000000000000
                ;mem[9895] <= 30'b000000001000000000000000010000
                ;mem[9896] <= 30'b000000001000000000000000100000
                ;mem[9897] <= 30'b000000001000000000000000110000
                ;mem[9898] <= 30'b000000001000000000000010010000
                ;mem[9899] <= 30'b000000001000000000000010100000
                ;mem[9900] <= 30'b000000001000000000000010110000
                ;mem[9901] <= 30'b000000001000000000000111000000
                ;mem[9902] <= 30'b000000001000000000000111010000
                ;mem[9903] <= 30'b000000001000000000001001100000
                ;mem[9904] <= 30'b000000001000000000001001110000
                ;mem[9905] <= 30'b000000001000000000001010000000
                ;mem[9906] <= 30'b000000001000000000010000110000
                ;mem[9907] <= 30'b000000001000000000010001000000
                ;mem[9908] <= 30'b000000001000000000011000000000
                ;mem[9909] <= 30'b000000001000000000011000010000
                ;mem[9910] <= 30'b000000001000000000011111000000
                ;mem[9911] <= 30'b000000001000000000011111010000
                ;mem[9912] <= 30'b000000001000000000100110000000
                ;mem[9913] <= 30'b000000001000000000100110010000
                ;mem[9914] <= 30'b000000001000000000101101000000
                ;mem[9915] <= 30'b000000001000000000101101010000
                ;mem[9916] <= 30'b000000001000000000110011110000
                ;mem[9917] <= 30'b000000001000000000110100000000
                ;mem[9918] <= 30'b000000001000000000111010110000
                ;mem[9919] <= 30'b000000001000000000111011000000
                ;mem[9920] <= 30'b000000010000000000000001000000
                ;mem[9921] <= 30'b000000010000000000000001010000
                ;mem[9922] <= 30'b000000010000000000000111110000
                ;mem[9923] <= 30'b000000010000000000001000000000
                ;mem[9924] <= 30'b000000010000000000001110110000
                ;mem[9925] <= 30'b000000010000000000001111000000
                ;mem[9926] <= 30'b000000010000000000010101110000
                ;mem[9927] <= 30'b000000010000000000010110000000
                ;mem[9928] <= 30'b000000010000000000011100100000
                ;mem[9929] <= 30'b000000010000000000011100110000
                ;mem[9930] <= 30'b000000010000000000100001010000
                ;mem[9931] <= 30'b000000010000000000100011010000
                ;mem[9932] <= 30'b000000010000000000100011100000
                ;mem[9933] <= 30'b000000010000000000100011110000
                ;mem[9934] <= 30'b000000010000000000100111110000
                ;mem[9935] <= 30'b000000010000000000101000000000
                ;mem[9936] <= 30'b000000010000000000101000010000
                ;mem[9937] <= 30'b000000010000000000101000100000
                ;mem[9938] <= 30'b000000010000000000101000110000
                ;mem[9939] <= 30'b000000010000000000101001000000
                ;mem[9940] <= 30'b000000010000000000101010010000
                ;mem[9941] <= 30'b000000010000000000101010100000
                ;mem[9942] <= 30'b000000010000000000101110100000
                ;mem[9943] <= 30'b000000010000000000101110110000
                ;mem[9944] <= 30'b000000010000000000101111000000
                ;mem[9945] <= 30'b000000010000000000101111100000
                ;mem[9946] <= 30'b000000010000000000101111110000
                ;mem[9947] <= 30'b000000010000000000110000000000
                ;mem[9948] <= 30'b000000010000000000110000010000
                ;mem[9949] <= 30'b000000010000000000110000100000
                ;mem[9950] <= 30'b000000010000000000110000110000
                ;mem[9951] <= 30'b000000010000000000110001000000
                ;mem[9952] <= 30'b000000010000000000110001010000
                ;mem[9953] <= 30'b000000010000000000110101100000
                ;mem[9954] <= 30'b000000010000000000110101110000
                ;mem[9955] <= 30'b000000010000000000110111010000
                ;mem[9956] <= 30'b000000010000000000110111100000
                ;mem[9957] <= 30'b000000010000000000110111110000
                ;mem[9958] <= 30'b000000010000000000111000000000
                ;mem[9959] <= 30'b000000010000000000111000010000
                ;mem[9960] <= 30'b000000010000000000111100100000
                ;mem[9961] <= 30'b000000010000000000111100110000
                ;mem[9962] <= 30'b000000010000000000111110000000
                ;mem[9963] <= 30'b000000010000000000111110010000
                ;mem[9964] <= 30'b000000010000000000111110100000
                ;mem[9965] <= 30'b000000010000000000111110110000
                ;mem[9966] <= 30'b000000010000000000111111000000
                ;mem[9967] <= 30'b000000010000000000111111010000
                ;mem[9968] <= 30'b000000010000000000111111100000
                ;mem[9969] <= 30'b000000000000000001000010100000
                ;mem[9970] <= 30'b000000000000000001000010110000
                ;mem[9971] <= 30'b000000000000000001000011000000
                ;mem[9972] <= 30'b000000000000000001000011100000
                ;mem[9973] <= 30'b000000000000000001000011110000
                ;mem[9974] <= 30'b000000000000000001000100000000
                ;mem[9975] <= 30'b000000000000000001000100010000
                ;mem[9976] <= 30'b000000000000000001000100100000
                ;mem[9977] <= 30'b000000000000000001000100110000
                ;mem[9978] <= 30'b000000000000000001000101000000
                ;mem[9979] <= 30'b000000000000000001000101010000
                ;mem[9980] <= 30'b000000000000000001001001100000
                ;mem[9981] <= 30'b000000000000000001001001110000
                ;mem[9982] <= 30'b000000000000000001001011010000
                ;mem[9983] <= 30'b000000000000000001001011100000
                ;mem[9984] <= 30'b000000000000000001001011110000
                ;mem[9985] <= 30'b000000000000000001001100000000
                ;mem[9986] <= 30'b000000000000000001001100010000
                ;mem[9987] <= 30'b000000000000000001010000100000
                ;mem[9988] <= 30'b000000000000000001010000110000
                ;mem[9989] <= 30'b000000000000000001010010000000
                ;mem[9990] <= 30'b000000000000000001010010010000
                ;mem[9991] <= 30'b000000000000000001010010100000
                ;mem[9992] <= 30'b000000000000000001010010110000
                ;mem[9993] <= 30'b000000000000000001010011000000
                ;mem[9994] <= 30'b000000000000000001010011010000
                ;mem[9995] <= 30'b000000000000000001010011100000
                ;mem[9996] <= 30'b000000000000000001010111100000
                ;mem[9997] <= 30'b000000000000000001010111110000
                ;mem[9998] <= 30'b000000000000000001011000000000
                ;mem[9999] <= 30'b000000000000000001011000010000
                ;mem[10000] <= 30'b000000000000000001011000100000
                ;mem[10001] <= 30'b000000000000000001011000110000
                ;mem[10002] <= 30'b000000000000000001011001000000
                ;mem[10003] <= 30'b000000000000000001011001010000
                ;mem[10004] <= 30'b000000000000000001011001100000
                ;mem[10005] <= 30'b000000000000000001011010010000
                ;mem[10006] <= 30'b000000000000000001011010100000
                ;mem[10007] <= 30'b000000000000000001011010110000
                ;mem[10008] <= 30'b000000000000000001011111000000
                ;mem[10009] <= 30'b000000000000000001011111010000
                ;mem[10010] <= 30'b000000000000000001011111100000
                ;mem[10011] <= 30'b000000000000000001011111110000
                ;mem[10012] <= 30'b000000000000000001100000000000
                ;mem[10013] <= 30'b000000000000000001100001100000
                ;mem[10014] <= 30'b000000000000000001100001110000
                ;mem[10015] <= 30'b000000000000000000101101010000
                ;mem[10016] <= 30'b000000000000000000101101100000
                ;mem[10017] <= 30'b000000000000000000101101110000
                ;mem[10018] <= 30'b000000000000000000101110000000
                ;mem[10019] <= 30'b000000000000000000101110010000
                ;mem[10020] <= 30'b000000000000000000101110100000
                ;mem[10021] <= 30'b000000000000000000101110110000
                ;mem[10022] <= 30'b000000000000000000110100000000
                ;mem[10023] <= 30'b000000000000000000110100010000
                ;mem[10024] <= 30'b000000000000000000110100100000
                ;mem[10025] <= 30'b000000000000000000110100110000
                ;mem[10026] <= 30'b000000000000000000110101000000
                ;mem[10027] <= 30'b000000000000000000110101010000
                ;mem[10028] <= 30'b000000000000000000110101100000
                ;mem[10029] <= 30'b000000000000000000110101110000
                ;mem[10030] <= 30'b000000000000000000111010110000
                ;mem[10031] <= 30'b000000000000000000111011000000
                ;mem[10032] <= 30'b000000000000000000111011010000
                ;mem[10033] <= 30'b000000000000000000111011100000
                ;mem[10034] <= 30'b000000000000000000111011110000
                ;mem[10035] <= 30'b000000000000000000111100000000
                ;mem[10036] <= 30'b000000000000000000111100010000
                ;mem[10037] <= 30'b000000000000000000111100100000
                ;mem[10038] <= 30'b000000000000000000111100110000
                ;mem[10039] <= 30'b000000001000000000000001010000
                ;mem[10040] <= 30'b000000001000000000000001100000
                ;mem[10041] <= 30'b000000001000000000000001110000
                ;mem[10042] <= 30'b000000001000000000000010000000
                ;mem[10043] <= 30'b000000001000000000000010010000
                ;mem[10044] <= 30'b000000001000000000000010100000
                ;mem[10045] <= 30'b000000001000000000000010110000
                ;mem[10046] <= 30'b000000001000000000001000000000
                ;mem[10047] <= 30'b000000001000000000001000010000
                ;mem[10048] <= 30'b000000001000000000001000100000
                ;mem[10049] <= 30'b000000001000000000001000110000
                ;mem[10050] <= 30'b000000001000000000001001000000
                ;mem[10051] <= 30'b000000001000000000001001010000
                ;mem[10052] <= 30'b000000001000000000001001100000
                ;mem[10053] <= 30'b000000001000000000001001110000
                ;mem[10054] <= 30'b000000001000000000001110110000
                ;mem[10055] <= 30'b000000001000000000001111000000
                ;mem[10056] <= 30'b000000001000000000001111010000
                ;mem[10057] <= 30'b000000001000000000001111100000
                ;mem[10058] <= 30'b000000001000000000001111110000
                ;mem[10059] <= 30'b000000001000000000010000000000
                ;mem[10060] <= 30'b000000001000000000010000010000
                ;mem[10061] <= 30'b000000001000000000010000100000
                ;mem[10062] <= 30'b000000001000000000010000110000
                ;mem[10063] <= 30'b000000001000000000010101110000
                ;mem[10064] <= 30'b000000001000000000010110000000
                ;mem[10065] <= 30'b000000001000000000010110010000
                ;mem[10066] <= 30'b000000001000000000010110100000
                ;mem[10067] <= 30'b000000001000000000010111010000
                ;mem[10068] <= 30'b000000001000000000010111100000
                ;mem[10069] <= 30'b000000001000000000010111110000
                ;mem[10070] <= 30'b000000001000000000011000000000
                ;mem[10071] <= 30'b000000001000000000011100100000
                ;mem[10072] <= 30'b000000001000000000011100110000
                ;mem[10073] <= 30'b000000001000000000011101000000
                ;mem[10074] <= 30'b000000001000000000011101010000
                ;mem[10075] <= 30'b000000001000000000011110010000
                ;mem[10076] <= 30'b000000001000000000011110100000
                ;mem[10077] <= 30'b000000001000000000011110110000
                ;mem[10078] <= 30'b000000001000000000011111000000
                ;mem[10079] <= 30'b000000001000000000100011110000
                ;mem[10080] <= 30'b000000001000000000100100000000
                ;mem[10081] <= 30'b000000001000000000100100010000
                ;mem[10082] <= 30'b000000001000000000100100110000
                ;mem[10083] <= 30'b000000001000000000100101000000
                ;mem[10084] <= 30'b000000001000000000100101010000
                ;mem[10085] <= 30'b000000001000000000100101100000
                ;mem[10086] <= 30'b000000001000000000100101110000
                ;mem[10087] <= 30'b000000001000000000101010110000
                ;mem[10088] <= 30'b000000001000000000101011000000
                ;mem[10089] <= 30'b000000001000000000101011010000
                ;mem[10090] <= 30'b000000001000000000101011100000
                ;mem[10091] <= 30'b000000001000000000101011110000
                ;mem[10092] <= 30'b000000001000000000101100000000
                ;mem[10093] <= 30'b000000001000000000101100010000
                ;mem[10094] <= 30'b000000001000000000101100100000
                ;mem[10095] <= 30'b000000001000000000101100110000
                ;mem[10096] <= 30'b000000001000000000110010010000
                ;mem[10097] <= 30'b000000001000000000110010100000
                ;mem[10098] <= 30'b000000001000000000110010110000
                ;mem[10099] <= 30'b000000001000000000110011000000
                ;mem[10100] <= 30'b000000001000000000110011010000
                ;mem[10101] <= 30'b000000001000000000110011100000
                ;mem[10102] <= 30'b000000001000000000110011110000
                ;mem[10103] <= 30'b000000001000000000111001100000
                ;mem[10104] <= 30'b000000001000000000111001110000
                ;mem[10105] <= 30'b000000001000000000111010000000
                ;mem[10106] <= 30'b000000001000000000111010010000
                ;mem[10107] <= 30'b000000001000000000111010100000
                ;mem[10108] <= 30'b000000010000000000000000000000
                ;mem[10109] <= 30'b000000010000000000000000010000
                ;mem[10110] <= 30'b000000010000000000000000100000
                ;mem[10111] <= 30'b000000010000000000000000110000
                ;mem[10112] <= 30'b000000010000000000000110010000
                ;mem[10113] <= 30'b000000010000000000000110100000
                ;mem[10114] <= 30'b000000010000000000000110110000
                ;mem[10115] <= 30'b000000010000000000000111000000
                ;mem[10116] <= 30'b000000010000000000000111010000
                ;mem[10117] <= 30'b000000010000000000000111100000
                ;mem[10118] <= 30'b000000010000000000000111110000
                ;mem[10119] <= 30'b000000010000000000001101100000
                ;mem[10120] <= 30'b000000010000000000001101110000
                ;mem[10121] <= 30'b000000010000000000001110000000
                ;mem[10122] <= 30'b000000010000000000001110010000
                ;mem[10123] <= 30'b000000010000000000001110100000
                ;mem[10124] <= 30'b000000010000000000010100100000
                ;mem[10125] <= 30'b000000010000000000010100110000
                ;mem[10126] <= 30'b000000010000000000010101000000
                ;mem[10127] <= 30'b000000010000000000010101010000
                ;mem[10128] <= 30'b000000010000000000011011010000
                ;mem[10129] <= 30'b000000010000000000011011100000
                ;mem[10130] <= 30'b000000010000000000011011110000
                ;mem[10131] <= 30'b000000010000000000011100000000
                ;mem[10132] <= 30'b000000010000000000011100010000
                ;mem[10133] <= 30'b000000010000000000100010000000
                ;mem[10134] <= 30'b000000010000000000100010010000
                ;mem[10135] <= 30'b000000010000000000100010100000
                ;mem[10136] <= 30'b000000010000000000100010110000
                ;mem[10137] <= 30'b000000010000000000101000110000
                ;mem[10138] <= 30'b000000010000000000101001000000
                ;mem[10139] <= 30'b000000010000000000101001010000
                ;mem[10140] <= 30'b000000010000000000101001100000
                ;mem[10141] <= 30'b000000010000000000101111100000
                ;mem[10142] <= 30'b000000010000000000101111110000
                ;mem[10143] <= 30'b000000010000000000110000000000
                ;mem[10144] <= 30'b000000010000000000110000010000
                ;mem[10145] <= 30'b000000010000000000110000100000
                ;mem[10146] <= 30'b000000010000000000110110010000
                ;mem[10147] <= 30'b000000010000000000110110100000
                ;mem[10148] <= 30'b000000010000000000110110110000
                ;mem[10149] <= 30'b000000010000000000110111000000
                ;mem[10150] <= 30'b000000010000000000110111010000
                ;mem[10151] <= 30'b000000010000000000111101000000
                ;mem[10152] <= 30'b000000010000000000111101010000
                ;mem[10153] <= 30'b000000010000000000111101100000
                ;mem[10154] <= 30'b000000010000000000111101110000
                ;mem[10155] <= 30'b000000010000000000111110000000
                ;mem[10156] <= 30'b000000000000000001000011100000
                ;mem[10157] <= 30'b000000000000000001000011110000
                ;mem[10158] <= 30'b000000000000000001000100000000
                ;mem[10159] <= 30'b000000000000000001000100010000
                ;mem[10160] <= 30'b000000000000000001000100100000
                ;mem[10161] <= 30'b000000000000000001001010010000
                ;mem[10162] <= 30'b000000000000000001001010100000
                ;mem[10163] <= 30'b000000000000000001001010110000
                ;mem[10164] <= 30'b000000000000000001001011000000
                ;mem[10165] <= 30'b000000000000000001001011010000
                ;mem[10166] <= 30'b000000000000000001010001000000
                ;mem[10167] <= 30'b000000000000000001010001010000
                ;mem[10168] <= 30'b000000000000000001010001100000
                ;mem[10169] <= 30'b000000000000000001010001110000
                ;mem[10170] <= 30'b000000000000000001010010000000
                ;mem[10171] <= 30'b000000000000000001011000000000
                ;mem[10172] <= 30'b000000000000000001011000010000
                ;mem[10173] <= 30'b000000000000000001011000100000
                ;mem[10174] <= 30'b000000000000000001011000110000
                ;mem[10175] <= 30'b000000000000000001011110110000
                ;mem[10176] <= 30'b000000000000000001011111000000
                ;mem[10177] <= 30'b000000000000000001011111010000
                ;mem[10178] <= 30'b000000000000000001011111100000
                ;mem[10179] <= 30'b000000000000000001011111110000
                ;mem[10180] <= 30'b000000000000000001100101110000
                ;mem[10181] <= 30'b000000000000000001100110000000
                ;mem[10182] <= 30'b000000000000000001100110010000
                ;mem[10183] <= 30'b000000000000000001100110100000
                ;mem[10184] <= 30'b000000000000000001101100110000
                ;mem[10185] <= 30'b000000000000000001101101000000
                ;mem[10186] <= 30'b000000000000000001101101010000
                ;mem[10187] <= 30'b000000000000000000100110010000
                ;mem[10188] <= 30'b000000000000000000100110100000
                ;mem[10189] <= 30'b000000000000000000101101010000
                ;mem[10190] <= 30'b000000000000000000101101100000
                ;mem[10191] <= 30'b000000000000000000101101110000
                ;mem[10192] <= 30'b000000000000000000110100010000
                ;mem[10193] <= 30'b000000000000000000110100100000
                ;mem[10194] <= 30'b000000000000000000110100110000
                ;mem[10195] <= 30'b000000000000000000111011000000
                ;mem[10196] <= 30'b000000000000000000111011010000
                ;mem[10197] <= 30'b000000000000000000111011100000
                ;mem[10198] <= 30'b000000000000000000111011110000
                ;mem[10199] <= 30'b000000001000000000000001010000
                ;mem[10200] <= 30'b000000001000000000000001100000
                ;mem[10201] <= 30'b000000001000000000000001110000
                ;mem[10202] <= 30'b000000001000000000001000010000
                ;mem[10203] <= 30'b000000001000000000001000100000
                ;mem[10204] <= 30'b000000001000000000001000110000
                ;mem[10205] <= 30'b000000001000000000001111000000
                ;mem[10206] <= 30'b000000001000000000001111010000
                ;mem[10207] <= 30'b000000001000000000001111100000
                ;mem[10208] <= 30'b000000001000000000001111110000
                ;mem[10209] <= 30'b000000001000000000010110000000
                ;mem[10210] <= 30'b000000001000000000010110010000
                ;mem[10211] <= 30'b000000001000000000010110100000
                ;mem[10212] <= 30'b000000001000000000010110110000
                ;mem[10213] <= 30'b000000001000000000011101000000
                ;mem[10214] <= 30'b000000001000000000011101010000
                ;mem[10215] <= 30'b000000001000000000011101100000
                ;mem[10216] <= 30'b000000001000000000011101110000
                ;mem[10217] <= 30'b000000001000000000100100000000
                ;mem[10218] <= 30'b000000001000000000100100010000
                ;mem[10219] <= 30'b000000001000000000100100100000
                ;mem[10220] <= 30'b000000001000000000100100110000
                ;mem[10221] <= 30'b000000001000000000101011000000
                ;mem[10222] <= 30'b000000001000000000101011010000
                ;mem[10223] <= 30'b000000001000000000101011100000
                ;mem[10224] <= 30'b000000001000000000101011110000
                ;mem[10225] <= 30'b000000001000000000110010010000
                ;mem[10226] <= 30'b000000001000000000110010100000
                ;mem[10227] <= 30'b000000001000000000110010110000
                ;mem[10228] <= 30'b000000001000000000111001010000
                ;mem[10229] <= 30'b000000001000000000111001100000
                ;mem[10230] <= 30'b000000001000000000111001110000
                ;mem[10231] <= 30'b000000010000000000000110010000
                ;mem[10232] <= 30'b000000010000000000000110100000
                ;mem[10233] <= 30'b000000010000000000000110110000
                ;mem[10234] <= 30'b000000010000000000001101010000
                ;mem[10235] <= 30'b000000010000000000001101100000
                ;mem[10236] <= 30'b000000010000000000001101110000
                ;mem[10237] <= 30'b000000010000000000010100010000
                ;mem[10238] <= 30'b000000010000000000010100100000
                ;mem[10239] <= 30'b000000010000000000010100110000
                ;mem[10240] <= 30'b000000010000000000011011010000
                ;mem[10241] <= 30'b000000010000000000011011100000
                ;mem[10242] <= 30'b000000010000000000011011110000
                ;mem[10243] <= 30'b000000010000000000100010010000
                ;mem[10244] <= 30'b000000010000000000100010100000
                ;mem[10245] <= 30'b000000010000000000100010110000
                ;mem[10246] <= 30'b000000010000000000101001010000
                ;mem[10247] <= 30'b000000010000000000101001100000
                ;mem[10248] <= 30'b000000010000000000101001110000
                ;mem[10249] <= 30'b000000010000000000110000010000
                ;mem[10250] <= 30'b000000010000000000110000100000
                ;mem[10251] <= 30'b000000010000000000110000110000
                ;mem[10252] <= 30'b000000010000000000110111010000
                ;mem[10253] <= 30'b000000010000000000110111100000
                ;mem[10254] <= 30'b000000010000000000110111110000
                ;mem[10255] <= 30'b000000010000000000111110000000
                ;mem[10256] <= 30'b000000010000000000111110010000
                ;mem[10257] <= 30'b000000010000000000111110100000
                ;mem[10258] <= 30'b000000000000000001000100010000
                ;mem[10259] <= 30'b000000000000000001000100100000
                ;mem[10260] <= 30'b000000000000000001000100110000
                ;mem[10261] <= 30'b000000000000000001001011010000
                ;mem[10262] <= 30'b000000000000000001001011100000
                ;mem[10263] <= 30'b000000000000000001001011110000
                ;mem[10264] <= 30'b000000000000000001010010000000
                ;mem[10265] <= 30'b000000000000000001010010010000
                ;mem[10266] <= 30'b000000000000000001010010100000
                ;mem[10267] <= 30'b000000000000000001011001000000
                ;mem[10268] <= 30'b000000000000000001011001010000
                ;mem[10269] <= 30'b000000000000000001011001100000
                ;mem[10270] <= 30'b000000000000000001100000000000
                ;mem[10271] <= 30'b000000000000000001100000010000
                ;mem[10272] <= 30'b000000000000000001100000100000
                ;mem[10273] <= 30'b000000000000000001100111010000
                ;mem[10274] <= 30'b000000000000000001100111100000
                ;mem[10275] <= 30'b000000000000000000110101100000
                ;mem[10276] <= 30'b000000000000000000110101110000
                ;mem[10277] <= 30'b000000000000000000111100010000
                ;mem[10278] <= 30'b000000000000000000111100100000
                ;mem[10279] <= 30'b000000000000000000111100110000
                ;mem[10280] <= 30'b000000001000000000001001100000
                ;mem[10281] <= 30'b000000001000000000001001110000
                ;mem[10282] <= 30'b000000001000000000010000010000
                ;mem[10283] <= 30'b000000001000000000010000100000
                ;mem[10284] <= 30'b000000001000000000010000110000
                ;mem[10285] <= 30'b000000001000000000010100000000
                ;mem[10286] <= 30'b000000001000000000010100010000
                ;mem[10287] <= 30'b000000001000000000010100100000
                ;mem[10288] <= 30'b000000001000000000010100110000
                ;mem[10289] <= 30'b000000001000000000010101010000
                ;mem[10290] <= 30'b000000001000000000010101100000
                ;mem[10291] <= 30'b000000001000000000010101110000
                ;mem[10292] <= 30'b000000001000000000010110000000
                ;mem[10293] <= 30'b000000001000000000010110010000
                ;mem[10294] <= 30'b000000001000000000010110100000
                ;mem[10295] <= 30'b000000001000000000010110110000
                ;mem[10296] <= 30'b000000001000000000010111000000
                ;mem[10297] <= 30'b000000001000000000010111010000
                ;mem[10298] <= 30'b000000001000000000010111100000
                ;mem[10299] <= 30'b000000001000000000010111110000
                ;mem[10300] <= 30'b000000001000000000011011010000
                ;mem[10301] <= 30'b000000001000000000011011100000
                ;mem[10302] <= 30'b000000001000000000011011110000
                ;mem[10303] <= 30'b000000001000000000011100000000
                ;mem[10304] <= 30'b000000001000000000011100010000
                ;mem[10305] <= 30'b000000001000000000011100100000
                ;mem[10306] <= 30'b000000001000000000011100110000
                ;mem[10307] <= 30'b000000001000000000011101000000
                ;mem[10308] <= 30'b000000001000000000011101010000
                ;mem[10309] <= 30'b000000001000000000011101100000
                ;mem[10310] <= 30'b000000001000000000011101110000
                ;mem[10311] <= 30'b000000001000000000011110000000
                ;mem[10312] <= 30'b000000001000000000011110010000
                ;mem[10313] <= 30'b000000001000000000011110100000
                ;mem[10314] <= 30'b000000001000000000100100110000
                ;mem[10315] <= 30'b000000001000000000100101000000
                ;mem[10316] <= 30'b000000001000000000100101010000
                ;mem[10317] <= 30'b000000001000000000101011110000
                ;mem[10318] <= 30'b000000001000000000101100000000
                ;mem[10319] <= 30'b000000001000000000110010110000
                ;mem[10320] <= 30'b000000001000000000110011000000
                ;mem[10321] <= 30'b000000001000000000111001100000
                ;mem[10322] <= 30'b000000001000000000111001110000
                ;mem[10323] <= 30'b000000001000000000111010000000
                ;mem[10324] <= 30'b000000010000000000000000000000
                ;mem[10325] <= 30'b000000010000000000000110110000
                ;mem[10326] <= 30'b000000010000000000000111000000
                ;mem[10327] <= 30'b000000010000000000001101100000
                ;mem[10328] <= 30'b000000010000000000001101110000
                ;mem[10329] <= 30'b000000010000000000001110000000
                ;mem[10330] <= 30'b000000010000000000010100100000
                ;mem[10331] <= 30'b000000010000000000010100110000
                ;mem[10332] <= 30'b000000010000000000010101000000
                ;mem[10333] <= 30'b000000010000000000010101010000
                ;mem[10334] <= 30'b000000010000000000010110000000
                ;mem[10335] <= 30'b000000010000000000011010100000
                ;mem[10336] <= 30'b000000010000000000011010110000
                ;mem[10337] <= 30'b000000010000000000011011000000
                ;mem[10338] <= 30'b000000010000000000011011010000
                ;mem[10339] <= 30'b000000010000000000011011100000
                ;mem[10340] <= 30'b000000010000000000011011110000
                ;mem[10341] <= 30'b000000010000000000011100000000
                ;mem[10342] <= 30'b000000010000000000011100010000
                ;mem[10343] <= 30'b000000010000000000011100100000
                ;mem[10344] <= 30'b000000010000000000011100110000
                ;mem[10345] <= 30'b000000010000000000011101000000
                ;mem[10346] <= 30'b000000010000000000100001110000
                ;mem[10347] <= 30'b000000010000000000100010000000
                ;mem[10348] <= 30'b000000010000000000100010010000
                ;mem[10349] <= 30'b000000010000000000100010100000
                ;mem[10350] <= 30'b000000010000000000100010110000
                ;mem[10351] <= 30'b000000010000000000100011000000
                ;mem[10352] <= 30'b000000010000000000100011010000
                ;mem[10353] <= 30'b000000010000000000100011100000
                ;mem[10354] <= 30'b000000010000000000101001100000
                ;mem[10355] <= 30'b000000010000000000101001110000
                ;mem[10356] <= 30'b000000010000000000110000100000
                ;mem[10357] <= 30'b000000010000000000110000110000
                ;mem[10358] <= 30'b000000010000000000110111100000
                ;mem[10359] <= 30'b000000010000000000110111110000
                ;mem[10360] <= 30'b000000010000000000111110010000
                ;mem[10361] <= 30'b000000010000000000111110100000
                ;mem[10362] <= 30'b000000010000000000111110110000
                ;mem[10363] <= 30'b000000000000000001000100100000
                ;mem[10364] <= 30'b000000000000000001000100110000
                ;mem[10365] <= 30'b000000000000000001001011100000
                ;mem[10366] <= 30'b000000000000000001001011110000
                ;mem[10367] <= 30'b000000000000000001010010010000
                ;mem[10368] <= 30'b000000000000000001010010100000
                ;mem[10369] <= 30'b000000000000000001010010110000
                ;mem[10370] <= 30'b000000000000000001011001010000
                ;mem[10371] <= 30'b000000000000000001011001100000
                ;mem[10372] <= 30'b000000000000000001011001110000
                ;mem[10373] <= 30'b000000000000000001100000010000
                ;mem[10374] <= 30'b000000000000000001100000100000
                ;mem[10375] <= 30'b000000000000000001100111010000
                ;mem[10376] <= 30'b000000000000000001100111100000
                ;mem[10377] <= 30'b000000000000000001101110010000
                ;mem[10378] <= 30'b000000000000000001101110100000
                ;mem[10379] <= 30'b000000000000000001110101100000
                ;mem[10380] <= 30'b000000000000000000011111010000
                ;mem[10381] <= 30'b000000000000000000011111100000
                ;mem[10382] <= 30'b000000000000000000011111110000
                ;mem[10383] <= 30'b000000000000000000100000000000
                ;mem[10384] <= 30'b000000000000000000100110000000
                ;mem[10385] <= 30'b000000000000000000100110010000
                ;mem[10386] <= 30'b000000000000000000100110100000
                ;mem[10387] <= 30'b000000000000000000100110110000
                ;mem[10388] <= 30'b000000000000000000100111000000
                ;mem[10389] <= 30'b000000000000000000101100110000
                ;mem[10390] <= 30'b000000000000000000101101000000
                ;mem[10391] <= 30'b000000000000000000101101110000
                ;mem[10392] <= 30'b000000000000000000101110000000
                ;mem[10393] <= 30'b000000000000000000101110010000
                ;mem[10394] <= 30'b000000000000000000110011100000
                ;mem[10395] <= 30'b000000000000000000110011110000
                ;mem[10396] <= 30'b000000000000000000110101000000
                ;mem[10397] <= 30'b000000000000000000111100000000
                ;mem[10398] <= 30'b000000001000000000000000110000
                ;mem[10399] <= 30'b000000001000000000000001000000
                ;mem[10400] <= 30'b000000001000000000000001110000
                ;mem[10401] <= 30'b000000001000000000000010000000
                ;mem[10402] <= 30'b000000001000000000000010010000
                ;mem[10403] <= 30'b000000001000000000000111100000
                ;mem[10404] <= 30'b000000001000000000000111110000
                ;mem[10405] <= 30'b000000001000000000001001000000
                ;mem[10406] <= 30'b000000001000000000010000000000
                ;mem[10407] <= 30'b000000001000000000010110110000
                ;mem[10408] <= 30'b000000001000000000010111000000
                ;mem[10409] <= 30'b000000001000000000011101100000
                ;mem[10410] <= 30'b000000001000000000011101110000
                ;mem[10411] <= 30'b000000001000000000011110000000
                ;mem[10412] <= 30'b000000001000000000100100010000
                ;mem[10413] <= 30'b000000001000000000100100100000
                ;mem[10414] <= 30'b000000001000000000100100110000
                ;mem[10415] <= 30'b000000001000000000101010110000
                ;mem[10416] <= 30'b000000001000000000101011000000
                ;mem[10417] <= 30'b000000001000000000101011010000
                ;mem[10418] <= 30'b000000001000000000101011100000
                ;mem[10419] <= 30'b000000001000000000110001100000
                ;mem[10420] <= 30'b000000001000000000110001110000
                ;mem[10421] <= 30'b000000001000000000110010000000
                ;mem[10422] <= 30'b000000001000000000110010010000
                ;mem[10423] <= 30'b000000001000000000110010100000
                ;mem[10424] <= 30'b000000001000000000110010110000
                ;mem[10425] <= 30'b000000001000000000111000110000
                ;mem[10426] <= 30'b000000001000000000111001000000
                ;mem[10427] <= 30'b000000001000000000111001010000
                ;mem[10428] <= 30'b000000001000000000111001100000
                ;mem[10429] <= 30'b000000001000000000111001110000
                ;mem[10430] <= 30'b000000001000000000111010000000
                ;mem[10431] <= 30'b000000010000000000000101100000
                ;mem[10432] <= 30'b000000010000000000000101110000
                ;mem[10433] <= 30'b000000010000000000000110000000
                ;mem[10434] <= 30'b000000010000000000000110010000
                ;mem[10435] <= 30'b000000010000000000000110100000
                ;mem[10436] <= 30'b000000010000000000000110110000
                ;mem[10437] <= 30'b000000010000000000001100110000
                ;mem[10438] <= 30'b000000010000000000001101000000
                ;mem[10439] <= 30'b000000010000000000001101010000
                ;mem[10440] <= 30'b000000010000000000001101100000
                ;mem[10441] <= 30'b000000010000000000001101110000
                ;mem[10442] <= 30'b000000010000000000001110000000
                ;mem[10443] <= 30'b000000010000000000010101000000
                ;mem[10444] <= 30'b000000010000000000010101010000
                ;mem[10445] <= 30'b000000010000000000010101100000
                ;mem[10446] <= 30'b000000010000000000011100010000
                ;mem[10447] <= 30'b000000010000000000011100100000
                ;mem[10448] <= 30'b000000010000000000011100110000
                ;mem[10449] <= 30'b000000010000000000100011100000
                ;mem[10450] <= 30'b000000010000000000100011110000
                ;mem[10451] <= 30'b000000010000000000101010100000
                ;mem[10452] <= 30'b000000010000000000101010110000
                ;mem[10453] <= 30'b000000010000000000110001100000
                ;mem[10454] <= 30'b000000010000000000110001110000
                ;mem[10455] <= 30'b000000010000000000111000010000
                ;mem[10456] <= 30'b000000010000000000111000100000
                ;mem[10457] <= 30'b000000010000000000111101000000
                ;mem[10458] <= 30'b000000010000000000111110110000
                ;mem[10459] <= 30'b000000010000000000111111000000
                ;mem[10460] <= 30'b000000010000000000111111010000
                ;mem[10461] <= 30'b000000010000000000111111100000
                ;mem[10462] <= 30'b000000000000000001000101100000
                ;mem[10463] <= 30'b000000000000000001000101110000
                ;mem[10464] <= 30'b000000000000000001001100010000
                ;mem[10465] <= 30'b000000000000000001001100100000
                ;mem[10466] <= 30'b000000000000000001010001000000
                ;mem[10467] <= 30'b000000000000000001010010110000
                ;mem[10468] <= 30'b000000000000000001010011000000
                ;mem[10469] <= 30'b000000000000000001010011010000
                ;mem[10470] <= 30'b000000000000000001010011100000
                ;mem[10471] <= 30'b000000000000000001011000000000
                ;mem[10472] <= 30'b000000000000000001011000010000
                ;mem[10473] <= 30'b000000000000000001011001100000
                ;mem[10474] <= 30'b000000000000000001011001110000
                ;mem[10475] <= 30'b000000000000000001011010000000
                ;mem[10476] <= 30'b000000000000000001011010010000
                ;mem[10477] <= 30'b000000000000000001011111000000
                ;mem[10478] <= 30'b000000000000000001011111010000
                ;mem[10479] <= 30'b000000000000000001011111100000
                ;mem[10480] <= 30'b000000000000000001011111110000
                ;mem[10481] <= 30'b000000000000000001100000000000
                ;mem[10482] <= 30'b000000000000000001100000010000
                ;mem[10483] <= 30'b000000000000000001100000100000
                ;mem[10484] <= 30'b000000000000000001100000110000
                ;mem[10485] <= 30'b000000000000000000110011110000
                ;mem[10486] <= 30'b000000000000000000110100000000
                ;mem[10487] <= 30'b000000000000000000110100010000
                ;mem[10488] <= 30'b000000000000000000110100100000
                ;mem[10489] <= 30'b000000000000000000111010010000
                ;mem[10490] <= 30'b000000000000000000111010100000
                ;mem[10491] <= 30'b000000000000000000111010110000
                ;mem[10492] <= 30'b000000000000000000111011000000
                ;mem[10493] <= 30'b000000000000000000111011010000
                ;mem[10494] <= 30'b000000000000000000111011100000
                ;mem[10495] <= 30'b000000000000000000111011110000
                ;mem[10496] <= 30'b000000000000000000111100000000
                ;mem[10497] <= 30'b000000001000000000000111110000
                ;mem[10498] <= 30'b000000001000000000001000000000
                ;mem[10499] <= 30'b000000001000000000001000010000
                ;mem[10500] <= 30'b000000001000000000001000100000
                ;mem[10501] <= 30'b000000001000000000001110010000
                ;mem[10502] <= 30'b000000001000000000001110100000
                ;mem[10503] <= 30'b000000001000000000001110110000
                ;mem[10504] <= 30'b000000001000000000001111000000
                ;mem[10505] <= 30'b000000001000000000001111010000
                ;mem[10506] <= 30'b000000001000000000001111100000
                ;mem[10507] <= 30'b000000001000000000001111110000
                ;mem[10508] <= 30'b000000001000000000010000000000
                ;mem[10509] <= 30'b000000001000000000010100110000
                ;mem[10510] <= 30'b000000001000000000010101000000
                ;mem[10511] <= 30'b000000001000000000010101010000
                ;mem[10512] <= 30'b000000001000000000010101100000
                ;mem[10513] <= 30'b000000001000000000010111000000
                ;mem[10514] <= 30'b000000001000000000010111010000
                ;mem[10515] <= 30'b000000001000000000010111100000
                ;mem[10516] <= 30'b000000001000000000011011100000
                ;mem[10517] <= 30'b000000001000000000011011110000
                ;mem[10518] <= 30'b000000001000000000011110010000
                ;mem[10519] <= 30'b000000001000000000011110100000
                ;mem[10520] <= 30'b000000001000000000100010010000
                ;mem[10521] <= 30'b000000001000000000100010100000
                ;mem[10522] <= 30'b000000001000000000100101010000
                ;mem[10523] <= 30'b000000001000000000100101100000
                ;mem[10524] <= 30'b000000001000000000101001010000
                ;mem[10525] <= 30'b000000001000000000101001100000
                ;mem[10526] <= 30'b000000001000000000101100010000
                ;mem[10527] <= 30'b000000001000000000101100100000
                ;mem[10528] <= 30'b000000001000000000110011010000
                ;mem[10529] <= 30'b000000001000000000110011100000
                ;mem[10530] <= 30'b000000001000000000111010010000
                ;mem[10531] <= 30'b000000001000000000111010100000
                ;mem[10532] <= 30'b000000010000000000000000010000
                ;mem[10533] <= 30'b000000010000000000000000100000
                ;mem[10534] <= 30'b000000010000000000000111010000
                ;mem[10535] <= 30'b000000010000000000000111100000
                ;mem[10536] <= 30'b000000010000000000001110010000
                ;mem[10537] <= 30'b000000010000000000001110100000
                ;mem[10538] <= 30'b000000010000000000010101000000
                ;mem[10539] <= 30'b000000010000000000010101010000
                ;mem[10540] <= 30'b000000010000000000011011110000
                ;mem[10541] <= 30'b000000010000000000011100000000
                ;mem[10542] <= 30'b000000010000000000100010100000
                ;mem[10543] <= 30'b000000010000000000100010110000
                ;mem[10544] <= 30'b000000010000000000101001000000
                ;mem[10545] <= 30'b000000010000000000101001010000
                ;mem[10546] <= 30'b000000010000000000101001100000
                ;mem[10547] <= 30'b000000010000000000101111110000
                ;mem[10548] <= 30'b000000010000000000110000000000
                ;mem[10549] <= 30'b000000010000000000110000010000
                ;mem[10550] <= 30'b000000010000000000110110100000
                ;mem[10551] <= 30'b000000010000000000110110110000
                ;mem[10552] <= 30'b000000010000000000110111000000
                ;mem[10553] <= 30'b000000010000000000110111010000
                ;mem[10554] <= 30'b000000010000000000110111100000
                ;mem[10555] <= 30'b000000010000000000110111110000
                ;mem[10556] <= 30'b000000010000000000111000000000
                ;mem[10557] <= 30'b000000010000000000111000010000
                ;mem[10558] <= 30'b000000010000000000111000100000
                ;mem[10559] <= 30'b000000010000000000111000110000
                ;mem[10560] <= 30'b000000010000000000111001000000
                ;mem[10561] <= 30'b000000010000000000111001010000
                ;mem[10562] <= 30'b000000010000000000111001100000
                ;mem[10563] <= 30'b000000010000000000111001110000
                ;mem[10564] <= 30'b000000010000000000111010000000
                ;mem[10565] <= 30'b000000010000000000111101100000
                ;mem[10566] <= 30'b000000010000000000111101110000
                ;mem[10567] <= 30'b000000010000000000111111010000
                ;mem[10568] <= 30'b000000010000000000111111100000
                ;mem[10569] <= 30'b000000010000000000111111110000
                ;mem[10570] <= 30'b000000000000000001000011110000
                ;mem[10571] <= 30'b000000000000000001000100000000
                ;mem[10572] <= 30'b000000000000000001000100010000
                ;mem[10573] <= 30'b000000000000000001001010100000
                ;mem[10574] <= 30'b000000000000000001001010110000
                ;mem[10575] <= 30'b000000000000000001001011000000
                ;mem[10576] <= 30'b000000000000000001001011010000
                ;mem[10577] <= 30'b000000000000000001001011100000
                ;mem[10578] <= 30'b000000000000000001001011110000
                ;mem[10579] <= 30'b000000000000000001001100000000
                ;mem[10580] <= 30'b000000000000000001001100010000
                ;mem[10581] <= 30'b000000000000000001001100100000
                ;mem[10582] <= 30'b000000000000000001001100110000
                ;mem[10583] <= 30'b000000000000000001001101000000
                ;mem[10584] <= 30'b000000000000000001001101010000
                ;mem[10585] <= 30'b000000000000000001001101100000
                ;mem[10586] <= 30'b000000000000000001001101110000
                ;mem[10587] <= 30'b000000000000000001001110000000
                ;mem[10588] <= 30'b000000000000000001010001100000
                ;mem[10589] <= 30'b000000000000000001010001110000
                ;mem[10590] <= 30'b000000000000000001010011010000
                ;mem[10591] <= 30'b000000000000000001010011100000
                ;mem[10592] <= 30'b000000000000000001010011110000
                ;mem[10593] <= 30'b000000000000000001010100010000
                ;mem[10594] <= 30'b000000000000000001010100100000
                ;mem[10595] <= 30'b000000000000000001010100110000
                ;mem[10596] <= 30'b000000000000000001010101000000
                ;mem[10597] <= 30'b000000000000000000101110000000
                ;mem[10598] <= 30'b000000000000000000101110010000
                ;mem[10599] <= 30'b000000000000000000110100110000
                ;mem[10600] <= 30'b000000000000000000110101000000
                ;mem[10601] <= 30'b000000000000000000110101010000
                ;mem[10602] <= 30'b000000000000000000110101100000
                ;mem[10603] <= 30'b000000000000000000111011100000
                ;mem[10604] <= 30'b000000000000000000111011110000
                ;mem[10605] <= 30'b000000000000000000111100000000
                ;mem[10606] <= 30'b000000000000000000111100010000
                ;mem[10607] <= 30'b000000000000000000111100100000
                ;mem[10608] <= 30'b000000001000000000000010000000
                ;mem[10609] <= 30'b000000001000000000000010010000
                ;mem[10610] <= 30'b000000001000000000001000110000
                ;mem[10611] <= 30'b000000001000000000001001000000
                ;mem[10612] <= 30'b000000001000000000001001010000
                ;mem[10613] <= 30'b000000001000000000001001100000
                ;mem[10614] <= 30'b000000001000000000001111100000
                ;mem[10615] <= 30'b000000001000000000001111110000
                ;mem[10616] <= 30'b000000001000000000010000000000
                ;mem[10617] <= 30'b000000001000000000010000010000
                ;mem[10618] <= 30'b000000001000000000010000100000
                ;mem[10619] <= 30'b000000001000000000010110010000
                ;mem[10620] <= 30'b000000001000000000010110100000
                ;mem[10621] <= 30'b000000001000000000010110110000
                ;mem[10622] <= 30'b000000001000000000010111100000
                ;mem[10623] <= 30'b000000001000000000011101000000
                ;mem[10624] <= 30'b000000001000000000011101010000
                ;mem[10625] <= 30'b000000001000000000011110100000
                ;mem[10626] <= 30'b000000001000000000011110110000
                ;mem[10627] <= 30'b000000001000000000100011110000
                ;mem[10628] <= 30'b000000001000000000100100000000
                ;mem[10629] <= 30'b000000001000000000100100010000
                ;mem[10630] <= 30'b000000001000000000100101010000
                ;mem[10631] <= 30'b000000001000000000100101100000
                ;mem[10632] <= 30'b000000001000000000100101110000
                ;mem[10633] <= 30'b000000001000000000101010100000
                ;mem[10634] <= 30'b000000001000000000101010110000
                ;mem[10635] <= 30'b000000001000000000101011000000
                ;mem[10636] <= 30'b000000001000000000101011100000
                ;mem[10637] <= 30'b000000001000000000101011110000
                ;mem[10638] <= 30'b000000001000000000101100000000
                ;mem[10639] <= 30'b000000001000000000101100010000
                ;mem[10640] <= 30'b000000001000000000101100100000
                ;mem[10641] <= 30'b000000001000000000110001100000
                ;mem[10642] <= 30'b000000001000000000110001110000
                ;mem[10643] <= 30'b000000001000000000110010000000
                ;mem[10644] <= 30'b000000001000000000110010010000
                ;mem[10645] <= 30'b000000001000000000110010100000
                ;mem[10646] <= 30'b000000001000000000110010110000
                ;mem[10647] <= 30'b000000001000000000110011000000
                ;mem[10648] <= 30'b000000001000000000110011010000
                ;mem[10649] <= 30'b000000001000000000110011100000
                ;mem[10650] <= 30'b000000001000000000111000100000
                ;mem[10651] <= 30'b000000001000000000111000110000
                ;mem[10652] <= 30'b000000001000000000111001000000
                ;mem[10653] <= 30'b000000001000000000111001010000
                ;mem[10654] <= 30'b000000001000000000111001100000
                ;mem[10655] <= 30'b000000001000000000111001110000
                ;mem[10656] <= 30'b000000001000000000111010000000
                ;mem[10657] <= 30'b000000001000000000111010010000
                ;mem[10658] <= 30'b000000010000000000000000000000
                ;mem[10659] <= 30'b000000010000000000000000010000
                ;mem[10660] <= 30'b000000010000000000000000100000
                ;mem[10661] <= 30'b000000010000000000000101100000
                ;mem[10662] <= 30'b000000010000000000000101110000
                ;mem[10663] <= 30'b000000010000000000000110000000
                ;mem[10664] <= 30'b000000010000000000000110010000
                ;mem[10665] <= 30'b000000010000000000000110100000
                ;mem[10666] <= 30'b000000010000000000000110110000
                ;mem[10667] <= 30'b000000010000000000000111000000
                ;mem[10668] <= 30'b000000010000000000000111010000
                ;mem[10669] <= 30'b000000010000000000000111100000
                ;mem[10670] <= 30'b000000010000000000001100100000
                ;mem[10671] <= 30'b000000010000000000001100110000
                ;mem[10672] <= 30'b000000010000000000001101000000
                ;mem[10673] <= 30'b000000010000000000001101010000
                ;mem[10674] <= 30'b000000010000000000001101100000
                ;mem[10675] <= 30'b000000010000000000001101110000
                ;mem[10676] <= 30'b000000010000000000001110000000
                ;mem[10677] <= 30'b000000010000000000001110010000
                ;mem[10678] <= 30'b000000010000000000010100100000
                ;mem[10679] <= 30'b000000010000000000010100110000
                ;mem[10680] <= 30'b000000010000000000010101000000
                ;mem[10681] <= 30'b000000010000000000011011010000
                ;mem[10682] <= 30'b000000010000000000011011100000
                ;mem[10683] <= 30'b000000010000000000011011110000
                ;mem[10684] <= 30'b000000010000000000100010010000
                ;mem[10685] <= 30'b000000010000000000100010100000
                ;mem[10686] <= 30'b000000010000000000101001000000
                ;mem[10687] <= 30'b000000010000000000101001010000
                ;mem[10688] <= 30'b000000010000000000101001100000
                ;mem[10689] <= 30'b000000010000000000110000000000
                ;mem[10690] <= 30'b000000010000000000110000010000
                ;mem[10691] <= 30'b000000010000000000110110110000
                ;mem[10692] <= 30'b000000010000000000110111000000
                ;mem[10693] <= 30'b000000010000000000110111010000
                ;mem[10694] <= 30'b000000010000000000111101110000
                ;mem[10695] <= 30'b000000010000000000111110000000
                ;mem[10696] <= 30'b000000000000000001000100000000
                ;mem[10697] <= 30'b000000000000000001000100010000
                ;mem[10698] <= 30'b000000000000000001001010110000
                ;mem[10699] <= 30'b000000000000000001001011000000
                ;mem[10700] <= 30'b000000000000000001001011010000
                ;mem[10701] <= 30'b000000000000000001010001110000
                ;mem[10702] <= 30'b000000000000000001010010000000
                ;mem[10703] <= 30'b000000000000000001011000110000
                ;mem[10704] <= 30'b000000000000000001011001000000
                ;mem[10705] <= 30'b000000000000000001011111110000
                ;mem[10706] <= 30'b000000000000000001100000000000
                ;mem[10707] <= 30'b000000000000000001100110110000
                ;mem[10708] <= 30'b000000000000000001100111000000
                ;mem[10709] <= 30'b000000000000000001100111010000
                ;mem[10710] <= 30'b000000000000000001100111100000
                ;mem[10711] <= 30'b000000000000000001101101110000
                ;mem[10712] <= 30'b000000000000000001101110000000
                ;mem[10713] <= 30'b000000000000000001101110010000
                ;mem[10714] <= 30'b000000000000000000110100110000
                ;mem[10715] <= 30'b000000000000000000110101000000
                ;mem[10716] <= 30'b000000000000000000110101010000
                ;mem[10717] <= 30'b000000000000000000110101100000
                ;mem[10718] <= 30'b000000000000000000110101110000
                ;mem[10719] <= 30'b000000000000000000110110000000
                ;mem[10720] <= 30'b000000000000000000110110010000
                ;mem[10721] <= 30'b000000000000000000111010010000
                ;mem[10722] <= 30'b000000000000000000111010100000
                ;mem[10723] <= 30'b000000000000000000111010110000
                ;mem[10724] <= 30'b000000000000000000111011000000
                ;mem[10725] <= 30'b000000000000000000111011010000
                ;mem[10726] <= 30'b000000000000000000111011100000
                ;mem[10727] <= 30'b000000000000000000111011110000
                ;mem[10728] <= 30'b000000000000000000111100000000
                ;mem[10729] <= 30'b000000000000000000111100010000
                ;mem[10730] <= 30'b000000000000000000111100100000
                ;mem[10731] <= 30'b000000000000000000111100110000
                ;mem[10732] <= 30'b000000000000000000111101000000
                ;mem[10733] <= 30'b000000000000000000111101010000
                ;mem[10734] <= 30'b000000001000000000001000110000
                ;mem[10735] <= 30'b000000001000000000001001000000
                ;mem[10736] <= 30'b000000001000000000001001010000
                ;mem[10737] <= 30'b000000001000000000001001100000
                ;mem[10738] <= 30'b000000001000000000001001110000
                ;mem[10739] <= 30'b000000001000000000001010000000
                ;mem[10740] <= 30'b000000001000000000001010010000
                ;mem[10741] <= 30'b000000001000000000001110010000
                ;mem[10742] <= 30'b000000001000000000001110100000
                ;mem[10743] <= 30'b000000001000000000001110110000
                ;mem[10744] <= 30'b000000001000000000001111000000
                ;mem[10745] <= 30'b000000001000000000001111010000
                ;mem[10746] <= 30'b000000001000000000001111100000
                ;mem[10747] <= 30'b000000001000000000001111110000
                ;mem[10748] <= 30'b000000001000000000010000000000
                ;mem[10749] <= 30'b000000001000000000010000010000
                ;mem[10750] <= 30'b000000001000000000010000100000
                ;mem[10751] <= 30'b000000001000000000010000110000
                ;mem[10752] <= 30'b000000001000000000010001000000
                ;mem[10753] <= 30'b000000001000000000010001010000
                ;mem[10754] <= 30'b000000001000000000010100100000
                ;mem[10755] <= 30'b000000001000000000010100110000
                ;mem[10756] <= 30'b000000001000000000010101000000
                ;mem[10757] <= 30'b000000001000000000010101010000
                ;mem[10758] <= 30'b000000001000000000010101100000
                ;mem[10759] <= 30'b000000001000000000010101110000
                ;mem[10760] <= 30'b000000001000000000010110000000
                ;mem[10761] <= 30'b000000001000000000010110010000
                ;mem[10762] <= 30'b000000001000000000010110100000
                ;mem[10763] <= 30'b000000001000000000010110110000
                ;mem[10764] <= 30'b000000001000000000010111000000
                ;mem[10765] <= 30'b000000001000000000010111010000
                ;mem[10766] <= 30'b000000001000000000010111100000
                ;mem[10767] <= 30'b000000001000000000010111110000
                ;mem[10768] <= 30'b000000001000000000011000000000
                ;mem[10769] <= 30'b000000001000000000011000010000
                ;mem[10770] <= 30'b000000001000000000011011100000
                ;mem[10771] <= 30'b000000001000000000011011110000
                ;mem[10772] <= 30'b000000001000000000011100000000
                ;mem[10773] <= 30'b000000001000000000011100010000
                ;mem[10774] <= 30'b000000001000000000011100100000
                ;mem[10775] <= 30'b000000001000000000011100110000
                ;mem[10776] <= 30'b000000001000000000011101000000
                ;mem[10777] <= 30'b000000001000000000011101010000
                ;mem[10778] <= 30'b000000001000000000011101100000
                ;mem[10779] <= 30'b000000001000000000011101110000
                ;mem[10780] <= 30'b000000001000000000011110000000
                ;mem[10781] <= 30'b000000001000000000011110010000
                ;mem[10782] <= 30'b000000001000000000011110100000
                ;mem[10783] <= 30'b000000001000000000011110110000
                ;mem[10784] <= 30'b000000001000000000011111000000
                ;mem[10785] <= 30'b000000001000000000011111010000
                ;mem[10786] <= 30'b000000001000000000100010100000
                ;mem[10787] <= 30'b000000001000000000100010110000
                ;mem[10788] <= 30'b000000001000000000100011000000
                ;mem[10789] <= 30'b000000001000000000100011010000
                ;mem[10790] <= 30'b000000001000000000100011100000
                ;mem[10791] <= 30'b000000001000000000100011110000
                ;mem[10792] <= 30'b000000001000000000100100000000
                ;mem[10793] <= 30'b000000001000000000100100010000
                ;mem[10794] <= 30'b000000001000000000100100100000
                ;mem[10795] <= 30'b000000001000000000100100110000
                ;mem[10796] <= 30'b000000001000000000100101000000
                ;mem[10797] <= 30'b000000001000000000100101010000
                ;mem[10798] <= 30'b000000001000000000100101100000
                ;mem[10799] <= 30'b000000001000000000100101110000
                ;mem[10800] <= 30'b000000001000000000100110000000
                ;mem[10801] <= 30'b000000001000000000100110010000
                ;mem[10802] <= 30'b000000001000000000101001110000
                ;mem[10803] <= 30'b000000001000000000101010000000
                ;mem[10804] <= 30'b000000001000000000101100010000
                ;mem[10805] <= 30'b000000001000000000101100100000
                ;mem[10806] <= 30'b000000001000000000101100110000
                ;mem[10807] <= 30'b000000001000000000101101000000
                ;mem[10808] <= 30'b000000001000000000101101010000
                ;mem[10809] <= 30'b000000001000000000110011000000
                ;mem[10810] <= 30'b000000001000000000110011010000
                ;mem[10811] <= 30'b000000001000000000110011100000
                ;mem[10812] <= 30'b000000001000000000110011110000
                ;mem[10813] <= 30'b000000001000000000110100000000
                ;mem[10814] <= 30'b000000001000000000110100010000
                ;mem[10815] <= 30'b000000001000000000111001110000
                ;mem[10816] <= 30'b000000001000000000111010000000
                ;mem[10817] <= 30'b000000001000000000111010010000
                ;mem[10818] <= 30'b000000001000000000111010100000
                ;mem[10819] <= 30'b000000001000000000111010110000
                ;mem[10820] <= 30'b000000001000000000111011000000
                ;mem[10821] <= 30'b000000010000000000000000010000
                ;mem[10822] <= 30'b000000010000000000000000100000
                ;mem[10823] <= 30'b000000010000000000000000110000
                ;mem[10824] <= 30'b000000010000000000000001000000
                ;mem[10825] <= 30'b000000010000000000000001010000
                ;mem[10826] <= 30'b000000010000000000000111000000
                ;mem[10827] <= 30'b000000010000000000000111010000
                ;mem[10828] <= 30'b000000010000000000000111100000
                ;mem[10829] <= 30'b000000010000000000000111110000
                ;mem[10830] <= 30'b000000010000000000001000000000
                ;mem[10831] <= 30'b000000010000000000001000010000
                ;mem[10832] <= 30'b000000010000000000001101110000
                ;mem[10833] <= 30'b000000010000000000001110000000
                ;mem[10834] <= 30'b000000010000000000001110010000
                ;mem[10835] <= 30'b000000010000000000001110100000
                ;mem[10836] <= 30'b000000010000000000001110110000
                ;mem[10837] <= 30'b000000010000000000001111000000
                ;mem[10838] <= 30'b000000010000000000010100100000
                ;mem[10839] <= 30'b000000010000000000010100110000
                ;mem[10840] <= 30'b000000010000000000010101000000
                ;mem[10841] <= 30'b000000010000000000010101010000
                ;mem[10842] <= 30'b000000010000000000010101100000
                ;mem[10843] <= 30'b000000010000000000010101110000
                ;mem[10844] <= 30'b000000010000000000011011010000
                ;mem[10845] <= 30'b000000010000000000011011100000
                ;mem[10846] <= 30'b000000010000000000011011110000
                ;mem[10847] <= 30'b000000010000000000011100000000
                ;mem[10848] <= 30'b000000010000000000011100010000
                ;mem[10849] <= 30'b000000010000000000011100100000
                ;mem[10850] <= 30'b000000010000000000011100110000
                ;mem[10851] <= 30'b000000010000000000100010000000
                ;mem[10852] <= 30'b000000010000000000100010010000
                ;mem[10853] <= 30'b000000010000000000100010100000
                ;mem[10854] <= 30'b000000010000000000100010110000
                ;mem[10855] <= 30'b000000010000000000100011000000
                ;mem[10856] <= 30'b000000010000000000100011010000
                ;mem[10857] <= 30'b000000010000000000101001000000
                ;mem[10858] <= 30'b000000010000000000101001010000
                ;mem[10859] <= 30'b000000010000000000101001100000
                ;mem[10860] <= 30'b000000010000000000101001110000
                ;mem[10861] <= 30'b000000010000000000101010000000
                ;mem[10862] <= 30'b000000010000000000101111100000
                ;mem[10863] <= 30'b000000010000000000101111110000
                ;mem[10864] <= 30'b000000010000000000110000000000
                ;mem[10865] <= 30'b000000010000000000110000010000
                ;mem[10866] <= 30'b000000010000000000110000100000
                ;mem[10867] <= 30'b000000010000000000110000110000
                ;mem[10868] <= 30'b000000010000000000110001000000
                ;mem[10869] <= 30'b000000010000000000110110100000
                ;mem[10870] <= 30'b000000010000000000110110110000
                ;mem[10871] <= 30'b000000010000000000110111000000
                ;mem[10872] <= 30'b000000010000000000110111010000
                ;mem[10873] <= 30'b000000010000000000110111100000
                ;mem[10874] <= 30'b000000010000000000111101010000
                ;mem[10875] <= 30'b000000010000000000111101100000
                ;mem[10876] <= 30'b000000010000000000111101110000
                ;mem[10877] <= 30'b000000010000000000111110000000
                ;mem[10878] <= 30'b000000010000000000111110010000
                ;mem[10879] <= 30'b000000010000000000111110100000
                ;mem[10880] <= 30'b000000000000000001000011100000
                ;mem[10881] <= 30'b000000000000000001000011110000
                ;mem[10882] <= 30'b000000000000000001000100000000
                ;mem[10883] <= 30'b000000000000000001000100010000
                ;mem[10884] <= 30'b000000000000000001000100100000
                ;mem[10885] <= 30'b000000000000000001000100110000
                ;mem[10886] <= 30'b000000000000000001000101000000
                ;mem[10887] <= 30'b000000000000000001001010100000
                ;mem[10888] <= 30'b000000000000000001001010110000
                ;mem[10889] <= 30'b000000000000000001001011000000
                ;mem[10890] <= 30'b000000000000000001001011010000
                ;mem[10891] <= 30'b000000000000000001001011100000
                ;mem[10892] <= 30'b000000000000000001010001010000
                ;mem[10893] <= 30'b000000000000000001010001100000
                ;mem[10894] <= 30'b000000000000000001010001110000
                ;mem[10895] <= 30'b000000000000000001010010000000
                ;mem[10896] <= 30'b000000000000000001010010010000
                ;mem[10897] <= 30'b000000000000000001010010100000
                ;mem[10898] <= 30'b000000000000000001011000000000
                ;mem[10899] <= 30'b000000000000000001011000010000
                ;mem[10900] <= 30'b000000000000000001011000100000
                ;mem[10901] <= 30'b000000000000000001011000110000
                ;mem[10902] <= 30'b000000000000000001011001000000
                ;mem[10903] <= 30'b000000000000000001011001010000
                ;mem[10904] <= 30'b000000000000000001011110110000
                ;mem[10905] <= 30'b000000000000000001011111000000
                ;mem[10906] <= 30'b000000000000000001011111010000
                ;mem[10907] <= 30'b000000000000000001011111100000
                ;mem[10908] <= 30'b000000000000000001011111110000
                ;mem[10909] <= 30'b000000000000000001100000000000
                ;mem[10910] <= 30'b000000000000000001100110000000
                ;mem[10911] <= 30'b000000000000000001100110010000
                ;mem[10912] <= 30'b000000000000000001100110100000
                ;mem[10913] <= 30'b000000000000000001100110110000
                ;mem[10914] <= 30'b000000000000000001100111000000
                ;mem[10915] <= 30'b000000000000000001101101000000
                ;mem[10916] <= 30'b000000000000000001101101010000
                ;mem[10917] <= 30'b000000000000000001101101100000
                ;mem[10918] <= 30'b000000000000000001101101110000
                ;mem[10919] <= 30'b000000000000000001110100100000
                ;mem[10920] <= 30'b000000000000000000110011100000
                ;mem[10921] <= 30'b000000000000000000110101000000
                ;mem[10922] <= 30'b000000000000000000111010010000
                ;mem[10923] <= 30'b000000000000000000111010100000
                ;mem[10924] <= 30'b000000000000000000111010110000
                ;mem[10925] <= 30'b000000000000000000111011000000
                ;mem[10926] <= 30'b000000000000000000111011010000
                ;mem[10927] <= 30'b000000000000000000111011100000
                ;mem[10928] <= 30'b000000000000000000111011110000
                ;mem[10929] <= 30'b000000000000000000111100000000
                ;mem[10930] <= 30'b000000000000000000111100010000
                ;mem[10931] <= 30'b000000001000000000000111100000
                ;mem[10932] <= 30'b000000001000000000001001000000
                ;mem[10933] <= 30'b000000001000000000001110010000
                ;mem[10934] <= 30'b000000001000000000001110100000
                ;mem[10935] <= 30'b000000001000000000001110110000
                ;mem[10936] <= 30'b000000001000000000001111000000
                ;mem[10937] <= 30'b000000001000000000001111010000
                ;mem[10938] <= 30'b000000001000000000001111100000
                ;mem[10939] <= 30'b000000001000000000001111110000
                ;mem[10940] <= 30'b000000001000000000010000000000
                ;mem[10941] <= 30'b000000001000000000010000010000
                ;mem[10942] <= 30'b000000001000000000010101010000
                ;mem[10943] <= 30'b000000001000000000010101100000
                ;mem[10944] <= 30'b000000001000000000010101110000
                ;mem[10945] <= 30'b000000001000000000010110000000
                ;mem[10946] <= 30'b000000001000000000010110010000
                ;mem[10947] <= 30'b000000001000000000010110100000
                ;mem[10948] <= 30'b000000001000000000010110110000
                ;mem[10949] <= 30'b000000001000000000010111000000
                ;mem[10950] <= 30'b000000001000000000010111010000
                ;mem[10951] <= 30'b000000001000000000011100010000
                ;mem[10952] <= 30'b000000001000000000011100100000
                ;mem[10953] <= 30'b000000001000000000011101000000
                ;mem[10954] <= 30'b000000001000000000011101010000
                ;mem[10955] <= 30'b000000001000000000011101100000
                ;mem[10956] <= 30'b000000001000000000011101110000
                ;mem[10957] <= 30'b000000001000000000011110000000
                ;mem[10958] <= 30'b000000001000000000011110010000
                ;mem[10959] <= 30'b000000001000000000100011010000
                ;mem[10960] <= 30'b000000001000000000100011100000
                ;mem[10961] <= 30'b000000001000000000100101000000
                ;mem[10962] <= 30'b000000001000000000100101010000
                ;mem[10963] <= 30'b000000001000000000101010010000
                ;mem[10964] <= 30'b000000001000000000101010100000
                ;mem[10965] <= 30'b000000001000000000101100000000
                ;mem[10966] <= 30'b000000001000000000101100010000
                ;mem[10967] <= 30'b000000001000000000110001010000
                ;mem[10968] <= 30'b000000001000000000110001100000
                ;mem[10969] <= 30'b000000001000000000110011000000
                ;mem[10970] <= 30'b000000001000000000110011010000
                ;mem[10971] <= 30'b000000001000000000110011100000
                ;mem[10972] <= 30'b000000001000000000111000010000
                ;mem[10973] <= 30'b000000001000000000111000100000
                ;mem[10974] <= 30'b000000001000000000111010000000
                ;mem[10975] <= 30'b000000001000000000111010010000
                ;mem[10976] <= 30'b000000001000000000111010100000
                ;mem[10977] <= 30'b000000001000000000111111010000
                ;mem[10978] <= 30'b000000001000000000111111100000
                ;mem[10979] <= 30'b000000010000000000000000000000
                ;mem[10980] <= 30'b000000010000000000000000010000
                ;mem[10981] <= 30'b000000010000000000000101010000
                ;mem[10982] <= 30'b000000010000000000000101100000
                ;mem[10983] <= 30'b000000010000000000000111000000
                ;mem[10984] <= 30'b000000010000000000000111010000
                ;mem[10985] <= 30'b000000010000000000000111100000
                ;mem[10986] <= 30'b000000010000000000001100010000
                ;mem[10987] <= 30'b000000010000000000001100100000
                ;mem[10988] <= 30'b000000010000000000001110000000
                ;mem[10989] <= 30'b000000010000000000001110010000
                ;mem[10990] <= 30'b000000010000000000001110100000
                ;mem[10991] <= 30'b000000010000000000010011010000
                ;mem[10992] <= 30'b000000010000000000010011100000
                ;mem[10993] <= 30'b000000010000000000010101000000
                ;mem[10994] <= 30'b000000010000000000010101010000
                ;mem[10995] <= 30'b000000010000000000010101100000
                ;mem[10996] <= 30'b000000010000000000011010100000
                ;mem[10997] <= 30'b000000010000000000011100000000
                ;mem[10998] <= 30'b000000010000000000011100010000
                ;mem[10999] <= 30'b000000010000000000011100100000
                ;mem[11000] <= 30'b000000010000000000100011000000
                ;mem[11001] <= 30'b000000010000000000100011010000
                ;mem[11002] <= 30'b000000010000000000100011100000
                ;mem[11003] <= 30'b000000010000000000101010000000
                ;mem[11004] <= 30'b000000010000000000101010010000
                ;mem[11005] <= 30'b000000010000000000101010100000
                ;mem[11006] <= 30'b000000010000000000110001000000
                ;mem[11007] <= 30'b000000010000000000110001010000
                ;mem[11008] <= 30'b000000010000000000110001100000
                ;mem[11009] <= 30'b000000010000000000111000000000
                ;mem[11010] <= 30'b000000010000000000111000010000
                ;mem[11011] <= 30'b000000010000000000111000100000
                ;mem[11012] <= 30'b000000010000000000111111000000
                ;mem[11013] <= 30'b000000010000000000111111010000
                ;mem[11014] <= 30'b000000010000000000111111100000
                ;mem[11015] <= 30'b000000000000000001000101000000
                ;mem[11016] <= 30'b000000000000000001000101010000
                ;mem[11017] <= 30'b000000000000000001000101100000
                ;mem[11018] <= 30'b000000000000000001001100000000
                ;mem[11019] <= 30'b000000000000000001001100010000
                ;mem[11020] <= 30'b000000000000000001001100100000
                ;mem[11021] <= 30'b000000000000000001010011000000
                ;mem[11022] <= 30'b000000000000000001010011010000
                ;mem[11023] <= 30'b000000000000000001010011100000
                ;mem[11024] <= 30'b000000000000000001011010000000
                ;mem[11025] <= 30'b000000000000000001011010010000
                ;mem[11026] <= 30'b000000000000000001011010100000
                ;mem[11027] <= 30'b000000000000000001100001000000
                ;mem[11028] <= 30'b000000000000000001100001010000
                ;mem[11029] <= 30'b000000000000000001100001100000
                ;mem[11030] <= 30'b000000000000000001101000000000
                ;mem[11031] <= 30'b000000000000000001101000010000
                ;mem[11032] <= 30'b000000000000000001101000100000
                ;mem[11033] <= 30'b000000000000000001101111000000
                ;mem[11034] <= 30'b000000000000000001101111010000
                ;mem[11035] <= 30'b000000000000000001101111100000
                ;mem[11036] <= 30'b000000000000000001110110010000
                ;mem[11037] <= 30'b000000000000000001110110100000
                ;mem[11038] <= 30'b000000000000000000011001000000
                ;mem[11039] <= 30'b000000000000000000011001010000
                ;mem[11040] <= 30'b000000000000000000011111100000
                ;mem[11041] <= 30'b000000000000000000011111110000
                ;mem[11042] <= 30'b000000000000000000100000000000
                ;mem[11043] <= 30'b000000000000000000100000010000
                ;mem[11044] <= 30'b000000000000000000100110010000
                ;mem[11045] <= 30'b000000000000000000100110100000
                ;mem[11046] <= 30'b000000000000000000100110110000
                ;mem[11047] <= 30'b000000000000000000100111000000
                ;mem[11048] <= 30'b000000000000000000100111010000
                ;mem[11049] <= 30'b000000000000000000101101000000
                ;mem[11050] <= 30'b000000000000000000101101010000
                ;mem[11051] <= 30'b000000000000000000101101100000
                ;mem[11052] <= 30'b000000000000000000101101110000
                ;mem[11053] <= 30'b000000000000000000101110000000
                ;mem[11054] <= 30'b000000000000000000101110010000
                ;mem[11055] <= 30'b000000000000000000110011110000
                ;mem[11056] <= 30'b000000000000000000110100000000
                ;mem[11057] <= 30'b000000000000000000110100010000
                ;mem[11058] <= 30'b000000000000000000110100100000
                ;mem[11059] <= 30'b000000000000000000111010100000
                ;mem[11060] <= 30'b000000000000000000111010110000
                ;mem[11061] <= 30'b000000000000000000111011000000
                ;mem[11062] <= 30'b000000000000000000111011010000
                ;mem[11063] <= 30'b000000001000000000000001000000
                ;mem[11064] <= 30'b000000001000000000000001010000
                ;mem[11065] <= 30'b000000001000000000000001100000
                ;mem[11066] <= 30'b000000001000000000000001110000
                ;mem[11067] <= 30'b000000001000000000000010000000
                ;mem[11068] <= 30'b000000001000000000000010010000
                ;mem[11069] <= 30'b000000001000000000000111110000
                ;mem[11070] <= 30'b000000001000000000001000000000
                ;mem[11071] <= 30'b000000001000000000001000010000
                ;mem[11072] <= 30'b000000001000000000001000100000
                ;mem[11073] <= 30'b000000001000000000001110100000
                ;mem[11074] <= 30'b000000001000000000001110110000
                ;mem[11075] <= 30'b000000001000000000001111000000
                ;mem[11076] <= 30'b000000001000000000001111010000
                ;mem[11077] <= 30'b000000001000000000010101100000
                ;mem[11078] <= 30'b000000001000000000010101110000
                ;mem[11079] <= 30'b000000001000000000010110000000
                ;mem[11080] <= 30'b000000001000000000011100010000
                ;mem[11081] <= 30'b000000001000000000011100100000
                ;mem[11082] <= 30'b000000001000000000011100110000
                ;mem[11083] <= 30'b000000001000000000100011010000
                ;mem[11084] <= 30'b000000001000000000100011100000
                ;mem[11085] <= 30'b000000001000000000100011110000
                ;mem[11086] <= 30'b000000001000000000101010010000
                ;mem[11087] <= 30'b000000001000000000101010100000
                ;mem[11088] <= 30'b000000001000000000101010110000
                ;mem[11089] <= 30'b000000001000000000110001010000
                ;mem[11090] <= 30'b000000001000000000110001100000
                ;mem[11091] <= 30'b000000001000000000110011100000
                ;mem[11092] <= 30'b000000001000000000110011110000
                ;mem[11093] <= 30'b000000001000000000111000010000
                ;mem[11094] <= 30'b000000001000000000111000100000
                ;mem[11095] <= 30'b000000001000000000111010000000
                ;mem[11096] <= 30'b000000001000000000111010010000
                ;mem[11097] <= 30'b000000001000000000111010100000
                ;mem[11098] <= 30'b000000001000000000111010110000
                ;mem[11099] <= 30'b000000001000000000111111010000
                ;mem[11100] <= 30'b000000001000000000111111100000
                ;mem[11101] <= 30'b000000010000000000000101010000
                ;mem[11102] <= 30'b000000010000000000000101100000
                ;mem[11103] <= 30'b000000010000000000000111100000
                ;mem[11104] <= 30'b000000010000000000000111110000
                ;mem[11105] <= 30'b000000010000000000001100010000
                ;mem[11106] <= 30'b000000010000000000001100100000
                ;mem[11107] <= 30'b000000010000000000001110000000
                ;mem[11108] <= 30'b000000010000000000001110010000
                ;mem[11109] <= 30'b000000010000000000001110100000
                ;mem[11110] <= 30'b000000010000000000001110110000
                ;mem[11111] <= 30'b000000010000000000010011010000
                ;mem[11112] <= 30'b000000010000000000010011100000
                ;mem[11113] <= 30'b000000010000000000010100110000
                ;mem[11114] <= 30'b000000010000000000010101000000
                ;mem[11115] <= 30'b000000010000000000010101010000
                ;mem[11116] <= 30'b000000010000000000010101100000
                ;mem[11117] <= 30'b000000010000000000010101110000
                ;mem[11118] <= 30'b000000010000000000010110000000
                ;mem[11119] <= 30'b000000010000000000011010010000
                ;mem[11120] <= 30'b000000010000000000011010100000
                ;mem[11121] <= 30'b000000010000000000011011110000
                ;mem[11122] <= 30'b000000010000000000011100000000
                ;mem[11123] <= 30'b000000010000000000011100010000
                ;mem[11124] <= 30'b000000010000000000011100100000
                ;mem[11125] <= 30'b000000010000000000011100110000
                ;mem[11126] <= 30'b000000010000000000011101000000
                ;mem[11127] <= 30'b000000010000000000100001010000
                ;mem[11128] <= 30'b000000010000000000100001100000
                ;mem[11129] <= 30'b000000010000000000100010100000
                ;mem[11130] <= 30'b000000010000000000100010110000
                ;mem[11131] <= 30'b000000010000000000100011000000
                ;mem[11132] <= 30'b000000010000000000100011110000
                ;mem[11133] <= 30'b000000010000000000100100000000
                ;mem[11134] <= 30'b000000010000000000101000010000
                ;mem[11135] <= 30'b000000010000000000101000100000
                ;mem[11136] <= 30'b000000010000000000101000110000
                ;mem[11137] <= 30'b000000010000000000101001100000
                ;mem[11138] <= 30'b000000010000000000101001110000
                ;mem[11139] <= 30'b000000010000000000101010110000
                ;mem[11140] <= 30'b000000010000000000101011000000
                ;mem[11141] <= 30'b000000010000000000101111100000
                ;mem[11142] <= 30'b000000010000000000101111110000
                ;mem[11143] <= 30'b000000010000000000110000000000
                ;mem[11144] <= 30'b000000010000000000110000100000
                ;mem[11145] <= 30'b000000010000000000110000110000
                ;mem[11146] <= 30'b000000010000000000110001000000
                ;mem[11147] <= 30'b000000010000000000110001100000
                ;mem[11148] <= 30'b000000010000000000110001110000
                ;mem[11149] <= 30'b000000010000000000110110100000
                ;mem[11150] <= 30'b000000010000000000110110110000
                ;mem[11151] <= 30'b000000010000000000110111000000
                ;mem[11152] <= 30'b000000010000000000110111010000
                ;mem[11153] <= 30'b000000010000000000110111100000
                ;mem[11154] <= 30'b000000010000000000110111110000
                ;mem[11155] <= 30'b000000010000000000111000000000
                ;mem[11156] <= 30'b000000010000000000111000010000
                ;mem[11157] <= 30'b000000010000000000111000100000
                ;mem[11158] <= 30'b000000010000000000111000110000
                ;mem[11159] <= 30'b000000010000000000111101110000
                ;mem[11160] <= 30'b000000010000000000111110000000
                ;mem[11161] <= 30'b000000010000000000111110010000
                ;mem[11162] <= 30'b000000010000000000111110100000
                ;mem[11163] <= 30'b000000010000000000111110110000
                ;mem[11164] <= 30'b000000010000000000111111000000
                ;mem[11165] <= 30'b000000010000000000111111010000
                ;mem[11166] <= 30'b000000010000000000111111100000
                ;mem[11167] <= 30'b000000000000000001000011100000
                ;mem[11168] <= 30'b000000000000000001000011110000
                ;mem[11169] <= 30'b000000000000000001000100000000
                ;mem[11170] <= 30'b000000000000000001000100100000
                ;mem[11171] <= 30'b000000000000000001000100110000
                ;mem[11172] <= 30'b000000000000000001000101000000
                ;mem[11173] <= 30'b000000000000000001000101100000
                ;mem[11174] <= 30'b000000000000000001000101110000
                ;mem[11175] <= 30'b000000000000000001001010100000
                ;mem[11176] <= 30'b000000000000000001001010110000
                ;mem[11177] <= 30'b000000000000000001001011000000
                ;mem[11178] <= 30'b000000000000000001001011010000
                ;mem[11179] <= 30'b000000000000000001001011100000
                ;mem[11180] <= 30'b000000000000000001001011110000
                ;mem[11181] <= 30'b000000000000000001001100000000
                ;mem[11182] <= 30'b000000000000000001001100010000
                ;mem[11183] <= 30'b000000000000000001001100100000
                ;mem[11184] <= 30'b000000000000000001001100110000
                ;mem[11185] <= 30'b000000000000000001010001110000
                ;mem[11186] <= 30'b000000000000000001010010000000
                ;mem[11187] <= 30'b000000000000000001010010010000
                ;mem[11188] <= 30'b000000000000000001010010100000
                ;mem[11189] <= 30'b000000000000000001010010110000
                ;mem[11190] <= 30'b000000000000000001010011000000
                ;mem[11191] <= 30'b000000000000000001010011010000
                ;mem[11192] <= 30'b000000000000000001010011100000
                ;mem[11193] <= 30'b000000000000000001011001010000
                ;mem[11194] <= 30'b000000000000000001011001100000
                ;mem[11195] <= 30'b000000000000000001011001110000
                ;mem[11196] <= 30'b000000000000000001011010000000
                ;mem[11197] <= 30'b000000000000000000011001000000
                ;mem[11198] <= 30'b000000000000000000011001010000
                ;mem[11199] <= 30'b000000000000000000011001100000
                ;mem[11200] <= 30'b000000000000000000011111000000
                ;mem[11201] <= 30'b000000000000000000011111010000
                ;mem[11202] <= 30'b000000000000000000011111100000
                ;mem[11203] <= 30'b000000000000000000011111110000
                ;mem[11204] <= 30'b000000000000000000100000000000
                ;mem[11205] <= 30'b000000000000000000100000010000
                ;mem[11206] <= 30'b000000000000000000100000100000
                ;mem[11207] <= 30'b000000000000000000100000110000
                ;mem[11208] <= 30'b000000000000000000100101010000
                ;mem[11209] <= 30'b000000000000000000100101100000
                ;mem[11210] <= 30'b000000000000000000100101110000
                ;mem[11211] <= 30'b000000000000000000100110000000
                ;mem[11212] <= 30'b000000000000000000100110010000
                ;mem[11213] <= 30'b000000000000000000100110100000
                ;mem[11214] <= 30'b000000000000000000100110110000
                ;mem[11215] <= 30'b000000000000000000100111000000
                ;mem[11216] <= 30'b000000000000000000100111010000
                ;mem[11217] <= 30'b000000000000000000100111100000
                ;mem[11218] <= 30'b000000000000000000100111110000
                ;mem[11219] <= 30'b000000000000000000101100000000
                ;mem[11220] <= 30'b000000000000000000101100010000
                ;mem[11221] <= 30'b000000000000000000101100100000
                ;mem[11222] <= 30'b000000000000000000101100110000
                ;mem[11223] <= 30'b000000000000000000101101000000
                ;mem[11224] <= 30'b000000000000000000101101010000
                ;mem[11225] <= 30'b000000000000000000101101100000
                ;mem[11226] <= 30'b000000000000000000101110010000
                ;mem[11227] <= 30'b000000000000000000101110100000
                ;mem[11228] <= 30'b000000000000000000101110110000
                ;mem[11229] <= 30'b000000000000000000110011010000
                ;mem[11230] <= 30'b000000000000000000110011100000
                ;mem[11231] <= 30'b000000000000000000110011110000
                ;mem[11232] <= 30'b000000000000000000110101100000
                ;mem[11233] <= 30'b000000000000000000110101110000
                ;mem[11234] <= 30'b000000000000000000111100100000
                ;mem[11235] <= 30'b000000000000000000111100110000
                ;mem[11236] <= 30'b000000001000000000000000000000
                ;mem[11237] <= 30'b000000001000000000000000010000
                ;mem[11238] <= 30'b000000001000000000000000100000
                ;mem[11239] <= 30'b000000001000000000000000110000
                ;mem[11240] <= 30'b000000001000000000000001000000
                ;mem[11241] <= 30'b000000001000000000000001010000
                ;mem[11242] <= 30'b000000001000000000000001100000
                ;mem[11243] <= 30'b000000001000000000000010010000
                ;mem[11244] <= 30'b000000001000000000000010100000
                ;mem[11245] <= 30'b000000001000000000000010110000
                ;mem[11246] <= 30'b000000001000000000000111010000
                ;mem[11247] <= 30'b000000001000000000000111100000
                ;mem[11248] <= 30'b000000001000000000000111110000
                ;mem[11249] <= 30'b000000001000000000001001100000
                ;mem[11250] <= 30'b000000001000000000001001110000
                ;mem[11251] <= 30'b000000001000000000010000100000
                ;mem[11252] <= 30'b000000001000000000010000110000
                ;mem[11253] <= 30'b000000001000000000010111100000
                ;mem[11254] <= 30'b000000001000000000010111110000
                ;mem[11255] <= 30'b000000001000000000011110100000
                ;mem[11256] <= 30'b000000001000000000011110110000
                ;mem[11257] <= 30'b000000001000000000100101010000
                ;mem[11258] <= 30'b000000001000000000100101100000
                ;mem[11259] <= 30'b000000001000000000100101110000
                ;mem[11260] <= 30'b000000001000000000101100010000
                ;mem[11261] <= 30'b000000001000000000101100100000
                ;mem[11262] <= 30'b000000001000000000101100110000
                ;mem[11263] <= 30'b000000001000000000110011000000
                ;mem[11264] <= 30'b000000001000000000110011010000
                ;mem[11265] <= 30'b000000001000000000110011100000
                ;mem[11266] <= 30'b000000001000000000111010000000
                ;mem[11267] <= 30'b000000001000000000111010010000
                ;mem[11268] <= 30'b000000001000000000111010100000
                ;mem[11269] <= 30'b000000010000000000000000010000
                ;mem[11270] <= 30'b000000010000000000000000100000
                ;mem[11271] <= 30'b000000010000000000000000110000
                ;mem[11272] <= 30'b000000010000000000000111000000
                ;mem[11273] <= 30'b000000010000000000000111010000
                ;mem[11274] <= 30'b000000010000000000000111100000
                ;mem[11275] <= 30'b000000010000000000001110000000
                ;mem[11276] <= 30'b000000010000000000001110010000
                ;mem[11277] <= 30'b000000010000000000001110100000
                ;mem[11278] <= 30'b000000010000000000010100110000
                ;mem[11279] <= 30'b000000010000000000010101000000
                ;mem[11280] <= 30'b000000010000000000010101010000
                ;mem[11281] <= 30'b000000010000000000010101100000
                ;mem[11282] <= 30'b000000010000000000011010010000
                ;mem[11283] <= 30'b000000010000000000011010100000
                ;mem[11284] <= 30'b000000010000000000011010110000
                ;mem[11285] <= 30'b000000010000000000011011000000
                ;mem[11286] <= 30'b000000010000000000011011010000
                ;mem[11287] <= 30'b000000010000000000011011100000
                ;mem[11288] <= 30'b000000010000000000011011110000
                ;mem[11289] <= 30'b000000010000000000011100000000
                ;mem[11290] <= 30'b000000010000000000011100010000
                ;mem[11291] <= 30'b000000010000000000100001000000
                ;mem[11292] <= 30'b000000010000000000100001010000
                ;mem[11293] <= 30'b000000010000000000100001100000
                ;mem[11294] <= 30'b000000010000000000100001110000
                ;mem[11295] <= 30'b000000010000000000100010000000
                ;mem[11296] <= 30'b000000010000000000100010010000
                ;mem[11297] <= 30'b000000010000000000100010100000
                ;mem[11298] <= 30'b000000010000000000100010110000
                ;mem[11299] <= 30'b000000010000000000100011000000
                ;mem[11300] <= 30'b000000010000000000100011010000
                ;mem[11301] <= 30'b000000010000000000100011100000
                ;mem[11302] <= 30'b000000010000000000100111110000
                ;mem[11303] <= 30'b000000010000000000101000000000
                ;mem[11304] <= 30'b000000010000000000101000010000
                ;mem[11305] <= 30'b000000010000000000101000100000
                ;mem[11306] <= 30'b000000010000000000101000110000
                ;mem[11307] <= 30'b000000010000000000101001000000
                ;mem[11308] <= 30'b000000010000000000101001010000
                ;mem[11309] <= 30'b000000010000000000101001100000
                ;mem[11310] <= 30'b000000010000000000101001110000
                ;mem[11311] <= 30'b000000010000000000101010000000
                ;mem[11312] <= 30'b000000010000000000101010010000
                ;mem[11313] <= 30'b000000010000000000101010100000
                ;mem[11314] <= 30'b000000010000000000101010110000
                ;mem[11315] <= 30'b000000010000000000101110100000
                ;mem[11316] <= 30'b000000010000000000101110110000
                ;mem[11317] <= 30'b000000010000000000101111000000
                ;mem[11318] <= 30'b000000010000000000101111010000
                ;mem[11319] <= 30'b000000010000000000101111100000
                ;mem[11320] <= 30'b000000010000000000101111110000
                ;mem[11321] <= 30'b000000010000000000110000000000
                ;mem[11322] <= 30'b000000010000000000110000010000
                ;mem[11323] <= 30'b000000010000000000110000100000
                ;mem[11324] <= 30'b000000010000000000110001000000
                ;mem[11325] <= 30'b000000010000000000110001010000
                ;mem[11326] <= 30'b000000010000000000110001100000
                ;mem[11327] <= 30'b000000010000000000110001110000
                ;mem[11328] <= 30'b000000010000000000110010000000
                ;mem[11329] <= 30'b000000010000000000110010010000
                ;mem[11330] <= 30'b000000010000000000110101100000
                ;mem[11331] <= 30'b000000010000000000110101110000
                ;mem[11332] <= 30'b000000010000000000110110000000
                ;mem[11333] <= 30'b000000010000000000110110010000
                ;mem[11334] <= 30'b000000010000000000110110100000
                ;mem[11335] <= 30'b000000010000000000110110110000
                ;mem[11336] <= 30'b000000010000000000110111000000
                ;mem[11337] <= 30'b000000010000000000110111010000
                ;mem[11338] <= 30'b000000010000000000111000110000
                ;mem[11339] <= 30'b000000010000000000111001000000
                ;mem[11340] <= 30'b000000010000000000111001010000
                ;mem[11341] <= 30'b000000010000000000111001100000
                ;mem[11342] <= 30'b000000010000000000111100100000
                ;mem[11343] <= 30'b000000010000000000111100110000
                ;mem[11344] <= 30'b000000010000000000111101000000
                ;mem[11345] <= 30'b000000010000000000111101010000
                ;mem[11346] <= 30'b000000010000000000111101100000
                ;mem[11347] <= 30'b000000010000000000111101110000
                ;mem[11348] <= 30'b000000000000000001000010100000
                ;mem[11349] <= 30'b000000000000000001000010110000
                ;mem[11350] <= 30'b000000000000000001000011000000
                ;mem[11351] <= 30'b000000000000000001000011010000
                ;mem[11352] <= 30'b000000000000000001000011100000
                ;mem[11353] <= 30'b000000000000000001000011110000
                ;mem[11354] <= 30'b000000000000000001000100000000
                ;mem[11355] <= 30'b000000000000000001000100010000
                ;mem[11356] <= 30'b000000000000000001000100100000
                ;mem[11357] <= 30'b000000000000000001000101000000
                ;mem[11358] <= 30'b000000000000000001000101010000
                ;mem[11359] <= 30'b000000000000000001000101100000
                ;mem[11360] <= 30'b000000000000000001000101110000
                ;mem[11361] <= 30'b000000000000000001000110000000
                ;mem[11362] <= 30'b000000000000000001000110010000
                ;mem[11363] <= 30'b000000000000000001001001100000
                ;mem[11364] <= 30'b000000000000000001001001110000
                ;mem[11365] <= 30'b000000000000000001001010000000
                ;mem[11366] <= 30'b000000000000000001001010010000
                ;mem[11367] <= 30'b000000000000000001001010100000
                ;mem[11368] <= 30'b000000000000000001001010110000
                ;mem[11369] <= 30'b000000000000000001001011000000
                ;mem[11370] <= 30'b000000000000000001001011010000
                ;mem[11371] <= 30'b000000000000000001001100110000
                ;mem[11372] <= 30'b000000000000000001001101000000
                ;mem[11373] <= 30'b000000000000000001001101010000
                ;mem[11374] <= 30'b000000000000000001001101100000
                ;mem[11375] <= 30'b000000000000000001010000100000
                ;mem[11376] <= 30'b000000000000000001010000110000
                ;mem[11377] <= 30'b000000000000000001010001000000
                ;mem[11378] <= 30'b000000000000000001010001010000
                ;mem[11379] <= 30'b000000000000000001010001100000
                ;mem[11380] <= 30'b000000000000000001010001110000
                ;mem[11381] <= 30'b000000000000000001010100010000
                ;mem[11382] <= 30'b000000000000000001010100100000
                ;mem[11383] <= 30'b000000000000000001010111110000
                ;mem[11384] <= 30'b000000000000000001011000000000
                ;mem[11385] <= 30'b000000000000000001011000010000
                ;mem[11386] <= 30'b000000000000000001011000100000
                ;mem[11387] <= 30'b000000000000000001011011100000
                ;mem[11388] <= 30'b000000000000000000110011010000
                ;mem[11389] <= 30'b000000000000000000111010000000
                ;mem[11390] <= 30'b000000000000000000111010010000
                ;mem[11391] <= 30'b000000000000000000111010100000
                ;mem[11392] <= 30'b000000000000000000111010110000
                ;mem[11393] <= 30'b000000000000000000111011000000
                ;mem[11394] <= 30'b000000000000000000111011010000
                ;mem[11395] <= 30'b000000000000000000111011100000
                ;mem[11396] <= 30'b000000000000000000111011110000
                ;mem[11397] <= 30'b000000000000000000111100000000
                ;mem[11398] <= 30'b000000000000000000111100010000
                ;mem[11399] <= 30'b000000000000000000111100100000
                ;mem[11400] <= 30'b000000001000000000000111010000
                ;mem[11401] <= 30'b000000001000000000001110000000
                ;mem[11402] <= 30'b000000001000000000001110010000
                ;mem[11403] <= 30'b000000001000000000001110100000
                ;mem[11404] <= 30'b000000001000000000001110110000
                ;mem[11405] <= 30'b000000001000000000001111000000
                ;mem[11406] <= 30'b000000001000000000001111010000
                ;mem[11407] <= 30'b000000001000000000001111100000
                ;mem[11408] <= 30'b000000001000000000001111110000
                ;mem[11409] <= 30'b000000001000000000010000000000
                ;mem[11410] <= 30'b000000001000000000010000010000
                ;mem[11411] <= 30'b000000001000000000010000100000
                ;mem[11412] <= 30'b000000001000000000010101010000
                ;mem[11413] <= 30'b000000001000000000010101100000
                ;mem[11414] <= 30'b000000001000000000010101110000
                ;mem[11415] <= 30'b000000001000000000010110000000
                ;mem[11416] <= 30'b000000001000000000010110010000
                ;mem[11417] <= 30'b000000001000000000010110100000
                ;mem[11418] <= 30'b000000001000000000010110110000
                ;mem[11419] <= 30'b000000001000000000010111000000
                ;mem[11420] <= 30'b000000001000000000010111010000
                ;mem[11421] <= 30'b000000001000000000010111100000
                ;mem[11422] <= 30'b000000001000000000010111110000
                ;mem[11423] <= 30'b000000001000000000011100000000
                ;mem[11424] <= 30'b000000001000000000011100010000
                ;mem[11425] <= 30'b000000001000000000011110010000
                ;mem[11426] <= 30'b000000001000000000011110100000
                ;mem[11427] <= 30'b000000001000000000011110110000
                ;mem[11428] <= 30'b000000001000000000100011000000
                ;mem[11429] <= 30'b000000001000000000100011010000
                ;mem[11430] <= 30'b000000001000000000100101010000
                ;mem[11431] <= 30'b000000001000000000100101100000
                ;mem[11432] <= 30'b000000001000000000101001110000
                ;mem[11433] <= 30'b000000001000000000101010000000
                ;mem[11434] <= 30'b000000001000000000101100010000
                ;mem[11435] <= 30'b000000001000000000101100100000
                ;mem[11436] <= 30'b000000001000000000110000110000
                ;mem[11437] <= 30'b000000001000000000110001000000
                ;mem[11438] <= 30'b000000001000000000110011010000
                ;mem[11439] <= 30'b000000001000000000110011100000
                ;mem[11440] <= 30'b000000001000000000111010000000
                ;mem[11441] <= 30'b000000001000000000111010010000
                ;mem[11442] <= 30'b000000001000000000111010100000
                ;mem[11443] <= 30'b000000010000000000000000010000
                ;mem[11444] <= 30'b000000010000000000000000100000
                ;mem[11445] <= 30'b000000010000000000000100110000
                ;mem[11446] <= 30'b000000010000000000000101000000
                ;mem[11447] <= 30'b000000010000000000000111010000
                ;mem[11448] <= 30'b000000010000000000000111100000
                ;mem[11449] <= 30'b000000010000000000001110000000
                ;mem[11450] <= 30'b000000010000000000001110010000
                ;mem[11451] <= 30'b000000010000000000001110100000
                ;mem[11452] <= 30'b000000010000000000010101000000
                ;mem[11453] <= 30'b000000010000000000010101010000
                ;mem[11454] <= 30'b000000010000000000010101100000
                ;mem[11455] <= 30'b000000010000000000011100000000
                ;mem[11456] <= 30'b000000010000000000011100010000
                ;mem[11457] <= 30'b000000010000000000100011000000
                ;mem[11458] <= 30'b000000010000000000100011010000
                ;mem[11459] <= 30'b000000010000000000101010000000
                ;mem[11460] <= 30'b000000010000000000101010010000
                ;mem[11461] <= 30'b000000010000000000110001000000
                ;mem[11462] <= 30'b000000010000000000110001010000
                ;mem[11463] <= 30'b000000010000000000111000000000
                ;mem[11464] <= 30'b000000010000000000111000010000
                ;mem[11465] <= 30'b000000010000000000111110110000
                ;mem[11466] <= 30'b000000010000000000111111000000
                ;mem[11467] <= 30'b000000010000000000111111010000
                ;mem[11468] <= 30'b000000000000000001000101000000
                ;mem[11469] <= 30'b000000000000000001000101010000
                ;mem[11470] <= 30'b000000000000000001001100000000
                ;mem[11471] <= 30'b000000000000000001001100010000
                ;mem[11472] <= 30'b000000000000000001010010110000
                ;mem[11473] <= 30'b000000000000000001010011000000
                ;mem[11474] <= 30'b000000000000000001010011010000
                ;mem[11475] <= 30'b000000000000000001011001110000
                ;mem[11476] <= 30'b000000000000000001011010000000
                ;mem[11477] <= 30'b000000000000000001011010010000
                ;mem[11478] <= 30'b000000000000000001100000110000
                ;mem[11479] <= 30'b000000000000000001100001000000
                ;mem[11480] <= 30'b000000000000000001100001010000
                ;mem[11481] <= 30'b000000000000000001100111110000
                ;mem[11482] <= 30'b000000000000000001101000000000
                ;mem[11483] <= 30'b000000000000000001101000010000
                ;mem[11484] <= 30'b000000000000000001101110110000
                ;mem[11485] <= 30'b000000000000000001101111000000
                ;mem[11486] <= 30'b000000000000000001110101110000
                ;mem[11487] <= 30'b000000000000000001110110000000
                ;mem[11488] <= 30'b000000000000000000101000000000
                ;mem[11489] <= 30'b000000000000000000101000010000
                ;mem[11490] <= 30'b000000000000000000101101110000
                ;mem[11491] <= 30'b000000000000000000101110000000
                ;mem[11492] <= 30'b000000000000000000101110110000
                ;mem[11493] <= 30'b000000000000000000101111000000
                ;mem[11494] <= 30'b000000000000000000101111010000
                ;mem[11495] <= 30'b000000000000000000101111100000
                ;mem[11496] <= 30'b000000000000000000110100010000
                ;mem[11497] <= 30'b000000000000000000110100100000
                ;mem[11498] <= 30'b000000000000000000110100110000
                ;mem[11499] <= 30'b000000000000000000110110000000
                ;mem[11500] <= 30'b000000000000000000110110010000
                ;mem[11501] <= 30'b000000000000000000110110100000
                ;mem[11502] <= 30'b000000000000000000111010100000
                ;mem[11503] <= 30'b000000000000000000111010110000
                ;mem[11504] <= 30'b000000000000000000111011000000
                ;mem[11505] <= 30'b000000000000000000111011010000
                ;mem[11506] <= 30'b000000000000000000111100110000
                ;mem[11507] <= 30'b000000000000000000111101000000
                ;mem[11508] <= 30'b000000000000000000111101010000
                ;mem[11509] <= 30'b000000001000000000000001110000
                ;mem[11510] <= 30'b000000001000000000000010000000
                ;mem[11511] <= 30'b000000001000000000000010110000
                ;mem[11512] <= 30'b000000001000000000000011000000
                ;mem[11513] <= 30'b000000001000000000000011010000
                ;mem[11514] <= 30'b000000001000000000000011100000
                ;mem[11515] <= 30'b000000001000000000001000010000
                ;mem[11516] <= 30'b000000001000000000001000100000
                ;mem[11517] <= 30'b000000001000000000001000110000
                ;mem[11518] <= 30'b000000001000000000001010000000
                ;mem[11519] <= 30'b000000001000000000001010010000
                ;mem[11520] <= 30'b000000001000000000001010100000
                ;mem[11521] <= 30'b000000001000000000001110100000
                ;mem[11522] <= 30'b000000001000000000001110110000
                ;mem[11523] <= 30'b000000001000000000001111000000
                ;mem[11524] <= 30'b000000001000000000001111010000
                ;mem[11525] <= 30'b000000001000000000010000110000
                ;mem[11526] <= 30'b000000001000000000010001000000
                ;mem[11527] <= 30'b000000001000000000010001010000
                ;mem[11528] <= 30'b000000001000000000010101000000
                ;mem[11529] <= 30'b000000001000000000010101010000
                ;mem[11530] <= 30'b000000001000000000010101100000
                ;mem[11531] <= 30'b000000001000000000010101110000
                ;mem[11532] <= 30'b000000001000000000010111010000
                ;mem[11533] <= 30'b000000001000000000010111100000
                ;mem[11534] <= 30'b000000001000000000010111110000
                ;mem[11535] <= 30'b000000001000000000011000000000
                ;mem[11536] <= 30'b000000001000000000011100000000
                ;mem[11537] <= 30'b000000001000000000011100010000
                ;mem[11538] <= 30'b000000001000000000011100100000
                ;mem[11539] <= 30'b000000001000000000011110000000
                ;mem[11540] <= 30'b000000001000000000011110010000
                ;mem[11541] <= 30'b000000001000000000011110100000
                ;mem[11542] <= 30'b000000001000000000100010110000
                ;mem[11543] <= 30'b000000001000000000100011000000
                ;mem[11544] <= 30'b000000001000000000100011010000
                ;mem[11545] <= 30'b000000001000000000100100110000
                ;mem[11546] <= 30'b000000001000000000100101000000
                ;mem[11547] <= 30'b000000001000000000100101010000
                ;mem[11548] <= 30'b000000001000000000101001110000
                ;mem[11549] <= 30'b000000001000000000101010000000
                ;mem[11550] <= 30'b000000001000000000101011100000
                ;mem[11551] <= 30'b000000001000000000101011110000
                ;mem[11552] <= 30'b000000001000000000101100000000
                ;mem[11553] <= 30'b000000001000000000110000110000
                ;mem[11554] <= 30'b000000001000000000110001000000
                ;mem[11555] <= 30'b000000001000000000110001010000
                ;mem[11556] <= 30'b000000001000000000110001100000
                ;mem[11557] <= 30'b000000001000000000110010010000
                ;mem[11558] <= 30'b000000001000000000110010100000
                ;mem[11559] <= 30'b000000001000000000110010110000
                ;mem[11560] <= 30'b000000001000000000111000000000
                ;mem[11561] <= 30'b000000001000000000111000010000
                ;mem[11562] <= 30'b000000001000000000111000100000
                ;mem[11563] <= 30'b000000001000000000111000110000
                ;mem[11564] <= 30'b000000001000000000111001000000
                ;mem[11565] <= 30'b000000001000000000111001010000
                ;mem[11566] <= 30'b000000001000000000111001100000
                ;mem[11567] <= 30'b000000001000000000111111100000
                ;mem[11568] <= 30'b000000001000000000111111110000
                ;mem[11569] <= 30'b000000010000000000000000000000
                ;mem[11570] <= 30'b000000010000000000000100110000
                ;mem[11571] <= 30'b000000010000000000000101000000
                ;mem[11572] <= 30'b000000010000000000000101010000
                ;mem[11573] <= 30'b000000010000000000000101100000
                ;mem[11574] <= 30'b000000010000000000000110010000
                ;mem[11575] <= 30'b000000010000000000000110100000
                ;mem[11576] <= 30'b000000010000000000000110110000
                ;mem[11577] <= 30'b000000010000000000001100000000
                ;mem[11578] <= 30'b000000010000000000001100010000
                ;mem[11579] <= 30'b000000010000000000001100100000
                ;mem[11580] <= 30'b000000010000000000001100110000
                ;mem[11581] <= 30'b000000010000000000001101000000
                ;mem[11582] <= 30'b000000010000000000001101010000
                ;mem[11583] <= 30'b000000010000000000001101100000
                ;mem[11584] <= 30'b000000010000000000010011100000
                ;mem[11585] <= 30'b000000010000000000010011110000
                ;mem[11586] <= 30'b000000010000000000010100000000
                ;mem[11587] <= 30'b000000010000000000010100010000
                ;mem[11588] <= 30'b000000010000000000010100100000
                ;mem[11589] <= 30'b000000010000000000010100110000
                ;mem[11590] <= 30'b000000010000000000011010110000
                ;mem[11591] <= 30'b000000010000000000011011000000
                ;mem[11592] <= 30'b000000010000000000011011010000
                ;mem[11593] <= 30'b000000010000000000011011100000
                ;mem[11594] <= 30'b000000010000000000011011110000
                ;mem[11595] <= 30'b000000010000000000011100000000
                ;mem[11596] <= 30'b000000010000000000011100010000
                ;mem[11597] <= 30'b000000010000000000100001110000
                ;mem[11598] <= 30'b000000010000000000100010000000
                ;mem[11599] <= 30'b000000010000000000100011010000
                ;mem[11600] <= 30'b000000010000000000100011100000
                ;mem[11601] <= 30'b000000010000000000100011110000
                ;mem[11602] <= 30'b000000010000000000101000110000
                ;mem[11603] <= 30'b000000010000000000101001000000
                ;mem[11604] <= 30'b000000010000000000101010100000
                ;mem[11605] <= 30'b000000010000000000101010110000
                ;mem[11606] <= 30'b000000010000000000101111110000
                ;mem[11607] <= 30'b000000010000000000110000000000
                ;mem[11608] <= 30'b000000010000000000110001110000
                ;mem[11609] <= 30'b000000010000000000110010000000
                ;mem[11610] <= 30'b000000010000000000110110110000
                ;mem[11611] <= 30'b000000010000000000110111000000
                ;mem[11612] <= 30'b000000010000000000111000100000
                ;mem[11613] <= 30'b000000010000000000111000110000
                ;mem[11614] <= 30'b000000010000000000111101110000
                ;mem[11615] <= 30'b000000010000000000111110000000
                ;mem[11616] <= 30'b000000010000000000111111100000
                ;mem[11617] <= 30'b000000010000000000111111110000
                ;mem[11618] <= 30'b000000000000000001000011110000
                ;mem[11619] <= 30'b000000000000000001000100000000
                ;mem[11620] <= 30'b000000000000000001000101110000
                ;mem[11621] <= 30'b000000000000000001000110000000
                ;mem[11622] <= 30'b000000000000000001001010110000
                ;mem[11623] <= 30'b000000000000000001001011000000
                ;mem[11624] <= 30'b000000000000000001001100100000
                ;mem[11625] <= 30'b000000000000000001001100110000
                ;mem[11626] <= 30'b000000000000000001010001110000
                ;mem[11627] <= 30'b000000000000000001010010000000
                ;mem[11628] <= 30'b000000000000000001010011100000
                ;mem[11629] <= 30'b000000000000000001010011110000
                ;mem[11630] <= 30'b000000000000000001011001000000
                ;mem[11631] <= 30'b000000000000000001011001010000
                ;mem[11632] <= 30'b000000000000000001011010100000
                ;mem[11633] <= 30'b000000000000000001011010110000
                ;mem[11634] <= 30'b000000000000000001100000010000
                ;mem[11635] <= 30'b000000000000000001100000100000
                ;mem[11636] <= 30'b000000000000000001100001000000
                ;mem[11637] <= 30'b000000000000000001100001010000
                ;mem[11638] <= 30'b000000000000000001100001100000
                ;mem[11639] <= 30'b000000000000000001100111100000
                ;mem[11640] <= 30'b000000000000000001100111110000
                ;mem[11641] <= 30'b000000000000000001101000000000
                ;mem[11642] <= 30'b000000000000000000100111110000
                ;mem[11643] <= 30'b000000000000000000101000000000
                ;mem[11644] <= 30'b000000000000000000101100000000
                ;mem[11645] <= 30'b000000000000000000101110100000
                ;mem[11646] <= 30'b000000000000000000101110110000
                ;mem[11647] <= 30'b000000000000000000101111000000
                ;mem[11648] <= 30'b000000000000000000101111010000
                ;mem[11649] <= 30'b000000000000000000110010110000
                ;mem[11650] <= 30'b000000000000000000110011000000
                ;mem[11651] <= 30'b000000000000000000110011010000
                ;mem[11652] <= 30'b000000000000000000110101100000
                ;mem[11653] <= 30'b000000000000000000110101110000
                ;mem[11654] <= 30'b000000000000000000110110000000
                ;mem[11655] <= 30'b000000000000000000110110010000
                ;mem[11656] <= 30'b000000000000000000111001110000
                ;mem[11657] <= 30'b000000000000000000111010000000
                ;mem[11658] <= 30'b000000000000000000111010010000
                ;mem[11659] <= 30'b000000000000000000111010100000
                ;mem[11660] <= 30'b000000000000000000111100100000
                ;mem[11661] <= 30'b000000000000000000111100110000
                ;mem[11662] <= 30'b000000000000000000111101000000
                ;mem[11663] <= 30'b000000000000000000111101010000
                ;mem[11664] <= 30'b000000001000000000000000000000
                ;mem[11665] <= 30'b000000001000000000000010100000
                ;mem[11666] <= 30'b000000001000000000000010110000
                ;mem[11667] <= 30'b000000001000000000000011000000
                ;mem[11668] <= 30'b000000001000000000000011010000
                ;mem[11669] <= 30'b000000001000000000000110110000
                ;mem[11670] <= 30'b000000001000000000000111000000
                ;mem[11671] <= 30'b000000001000000000000111010000
                ;mem[11672] <= 30'b000000001000000000001001100000
                ;mem[11673] <= 30'b000000001000000000001001110000
                ;mem[11674] <= 30'b000000001000000000001010000000
                ;mem[11675] <= 30'b000000001000000000001010010000
                ;mem[11676] <= 30'b000000001000000000001101110000
                ;mem[11677] <= 30'b000000001000000000001110000000
                ;mem[11678] <= 30'b000000001000000000001110010000
                ;mem[11679] <= 30'b000000001000000000001110100000
                ;mem[11680] <= 30'b000000001000000000010000100000
                ;mem[11681] <= 30'b000000001000000000010000110000
                ;mem[11682] <= 30'b000000001000000000010001000000
                ;mem[11683] <= 30'b000000001000000000010001010000
                ;mem[11684] <= 30'b000000001000000000010100110000
                ;mem[11685] <= 30'b000000001000000000010101000000
                ;mem[11686] <= 30'b000000001000000000010101010000
                ;mem[11687] <= 30'b000000001000000000010101100000
                ;mem[11688] <= 30'b000000001000000000010111010000
                ;mem[11689] <= 30'b000000001000000000010111100000
                ;mem[11690] <= 30'b000000001000000000010111110000
                ;mem[11691] <= 30'b000000001000000000011000000000
                ;mem[11692] <= 30'b000000001000000000011011110000
                ;mem[11693] <= 30'b000000001000000000011100000000
                ;mem[11694] <= 30'b000000001000000000011100010000
                ;mem[11695] <= 30'b000000001000000000011100100000
                ;mem[11696] <= 30'b000000001000000000011110010000
                ;mem[11697] <= 30'b000000001000000000011110100000
                ;mem[11698] <= 30'b000000001000000000011110110000
                ;mem[11699] <= 30'b000000001000000000011111000000
                ;mem[11700] <= 30'b000000001000000000100010100000
                ;mem[11701] <= 30'b000000001000000000100010110000
                ;mem[11702] <= 30'b000000001000000000100011000000
                ;mem[11703] <= 30'b000000001000000000100011010000
                ;mem[11704] <= 30'b000000001000000000100011100000
                ;mem[11705] <= 30'b000000001000000000100100110000
                ;mem[11706] <= 30'b000000001000000000100101000000
                ;mem[11707] <= 30'b000000001000000000100101010000
                ;mem[11708] <= 30'b000000001000000000100101100000
                ;mem[11709] <= 30'b000000001000000000100101110000
                ;mem[11710] <= 30'b000000001000000000100110000000
                ;mem[11711] <= 30'b000000001000000000101001100000
                ;mem[11712] <= 30'b000000001000000000101001110000
                ;mem[11713] <= 30'b000000001000000000101010000000
                ;mem[11714] <= 30'b000000001000000000101010010000
                ;mem[11715] <= 30'b000000001000000000101010100000
                ;mem[11716] <= 30'b000000001000000000101010110000
                ;mem[11717] <= 30'b000000001000000000101011000000
                ;mem[11718] <= 30'b000000001000000000101011010000
                ;mem[11719] <= 30'b000000001000000000101011100000
                ;mem[11720] <= 30'b000000001000000000101011110000
                ;mem[11721] <= 30'b000000001000000000101100000000
                ;mem[11722] <= 30'b000000001000000000101100010000
                ;mem[11723] <= 30'b000000001000000000101100100000
                ;mem[11724] <= 30'b000000001000000000101100110000
                ;mem[11725] <= 30'b000000001000000000110000100000
                ;mem[11726] <= 30'b000000001000000000110000110000
                ;mem[11727] <= 30'b000000001000000000110001000000
                ;mem[11728] <= 30'b000000001000000000110001010000
                ;mem[11729] <= 30'b000000001000000000110001100000
                ;mem[11730] <= 30'b000000001000000000110001110000
                ;mem[11731] <= 30'b000000001000000000110010000000
                ;mem[11732] <= 30'b000000001000000000110010010000
                ;mem[11733] <= 30'b000000001000000000110010100000
                ;mem[11734] <= 30'b000000001000000000110010110000
                ;mem[11735] <= 30'b000000001000000000110011000000
                ;mem[11736] <= 30'b000000001000000000110011010000
                ;mem[11737] <= 30'b000000001000000000110011100000
                ;mem[11738] <= 30'b000000001000000000110011110000
                ;mem[11739] <= 30'b000000001000000000110111100000
                ;mem[11740] <= 30'b000000001000000000110111110000
                ;mem[11741] <= 30'b000000001000000000111000000000
                ;mem[11742] <= 30'b000000001000000000111000010000
                ;mem[11743] <= 30'b000000001000000000111000100000
                ;mem[11744] <= 30'b000000001000000000111000110000
                ;mem[11745] <= 30'b000000001000000000111001000000
                ;mem[11746] <= 30'b000000001000000000111001010000
                ;mem[11747] <= 30'b000000001000000000111001100000
                ;mem[11748] <= 30'b000000001000000000111001110000
                ;mem[11749] <= 30'b000000001000000000111010000000
                ;mem[11750] <= 30'b000000001000000000111010010000
                ;mem[11751] <= 30'b000000001000000000111010100000
                ;mem[11752] <= 30'b000000001000000000111010110000
                ;mem[11753] <= 30'b000000001000000000111110100000
                ;mem[11754] <= 30'b000000001000000000111110110000
                ;mem[11755] <= 30'b000000001000000000111111000000
                ;mem[11756] <= 30'b000000001000000000111111010000
                ;mem[11757] <= 30'b000000001000000000111111100000
                ;mem[11758] <= 30'b000000001000000000111111110000
                ;mem[11759] <= 30'b000000010000000000000000000000
                ;mem[11760] <= 30'b000000010000000000000000010000
                ;mem[11761] <= 30'b000000010000000000000000100000
                ;mem[11762] <= 30'b000000010000000000000000110000
                ;mem[11763] <= 30'b000000010000000000000100100000
                ;mem[11764] <= 30'b000000010000000000000100110000
                ;mem[11765] <= 30'b000000010000000000000101000000
                ;mem[11766] <= 30'b000000010000000000000101010000
                ;mem[11767] <= 30'b000000010000000000000101100000
                ;mem[11768] <= 30'b000000010000000000000101110000
                ;mem[11769] <= 30'b000000010000000000000110000000
                ;mem[11770] <= 30'b000000010000000000000110010000
                ;mem[11771] <= 30'b000000010000000000000110100000
                ;mem[11772] <= 30'b000000010000000000000110110000
                ;mem[11773] <= 30'b000000010000000000000111000000
                ;mem[11774] <= 30'b000000010000000000000111010000
                ;mem[11775] <= 30'b000000010000000000000111100000
                ;mem[11776] <= 30'b000000010000000000000111110000
                ;mem[11777] <= 30'b000000010000000000001011100000
                ;mem[11778] <= 30'b000000010000000000001011110000
                ;mem[11779] <= 30'b000000010000000000001100000000
                ;mem[11780] <= 30'b000000010000000000001100010000
                ;mem[11781] <= 30'b000000010000000000001100100000
                ;mem[11782] <= 30'b000000010000000000001100110000
                ;mem[11783] <= 30'b000000010000000000001101000000
                ;mem[11784] <= 30'b000000010000000000001101010000
                ;mem[11785] <= 30'b000000010000000000001101100000
                ;mem[11786] <= 30'b000000010000000000001101110000
                ;mem[11787] <= 30'b000000010000000000001110000000
                ;mem[11788] <= 30'b000000010000000000001110010000
                ;mem[11789] <= 30'b000000010000000000001110100000
                ;mem[11790] <= 30'b000000010000000000001110110000
                ;mem[11791] <= 30'b000000010000000000010010100000
                ;mem[11792] <= 30'b000000010000000000010010110000
                ;mem[11793] <= 30'b000000010000000000010011000000
                ;mem[11794] <= 30'b000000010000000000010011010000
                ;mem[11795] <= 30'b000000010000000000010011100000
                ;mem[11796] <= 30'b000000010000000000010011110000
                ;mem[11797] <= 30'b000000010000000000010100000000
                ;mem[11798] <= 30'b000000010000000000010100010000
                ;mem[11799] <= 30'b000000010000000000010100100000
                ;mem[11800] <= 30'b000000010000000000010100110000
                ;mem[11801] <= 30'b000000010000000000010101000000
                ;mem[11802] <= 30'b000000010000000000010101010000
                ;mem[11803] <= 30'b000000010000000000010101100000
                ;mem[11804] <= 30'b000000010000000000011001110000
                ;mem[11805] <= 30'b000000010000000000011010000000
                ;mem[11806] <= 30'b000000010000000000011010010000
                ;mem[11807] <= 30'b000000010000000000011010100000
                ;mem[11808] <= 30'b000000010000000000011010110000
                ;mem[11809] <= 30'b000000010000000000011011000000
                ;mem[11810] <= 30'b000000010000000000011011010000
                ;mem[11811] <= 30'b000000010000000000011011110000
                ;mem[11812] <= 30'b000000010000000000011100000000
                ;mem[11813] <= 30'b000000010000000000011100010000
                ;mem[11814] <= 30'b000000010000000000011100100000
                ;mem[11815] <= 30'b000000010000000000100001000000
                ;mem[11816] <= 30'b000000010000000000100001010000
                ;mem[11817] <= 30'b000000010000000000100001100000
                ;mem[11818] <= 30'b000000010000000000100011000000
                ;mem[11819] <= 30'b000000010000000000100011010000
                ;mem[11820] <= 30'b000000010000000000100011100000
                ;mem[11821] <= 30'b000000010000000000100011110000
                ;mem[11822] <= 30'b000000010000000000100100000000
                ;mem[11823] <= 30'b000000010000000000101010000000
                ;mem[11824] <= 30'b000000010000000000101010010000
                ;mem[11825] <= 30'b000000010000000000101010100000
                ;mem[11826] <= 30'b000000010000000000101010110000
                ;mem[11827] <= 30'b000000010000000000101011000000
                ;mem[11828] <= 30'b000000010000000000110001000000
                ;mem[11829] <= 30'b000000010000000000110001010000
                ;mem[11830] <= 30'b000000010000000000110001100000
                ;mem[11831] <= 30'b000000010000000000110001110000
                ;mem[11832] <= 30'b000000010000000000110111110000
                ;mem[11833] <= 30'b000000010000000000111000000000
                ;mem[11834] <= 30'b000000010000000000111000010000
                ;mem[11835] <= 30'b000000010000000000111000100000
                ;mem[11836] <= 30'b000000010000000000111110110000
                ;mem[11837] <= 30'b000000010000000000111111000000
                ;mem[11838] <= 30'b000000010000000000111111010000
                ;mem[11839] <= 30'b000000010000000000111111100000
                ;mem[11840] <= 30'b000000000000000001000101000000
                ;mem[11841] <= 30'b000000000000000001000101010000
                ;mem[11842] <= 30'b000000000000000001000101100000
                ;mem[11843] <= 30'b000000000000000001000101110000
                ;mem[11844] <= 30'b000000000000000001001011110000
                ;mem[11845] <= 30'b000000000000000001001100000000
                ;mem[11846] <= 30'b000000000000000001001100010000
                ;mem[11847] <= 30'b000000000000000001001100100000
                ;mem[11848] <= 30'b000000000000000001010010110000
                ;mem[11849] <= 30'b000000000000000001010011000000
                ;mem[11850] <= 30'b000000000000000001010011010000
                ;mem[11851] <= 30'b000000000000000001010011100000
                ;mem[11852] <= 30'b000000000000000001011001110000
                ;mem[11853] <= 30'b000000000000000001011010000000
                ;mem[11854] <= 30'b000000000000000001011010010000
                ;mem[11855] <= 30'b000000000000000001100000110000
                ;mem[11856] <= 30'b000000000000000001100001000000
                ;mem[11857] <= 30'b000000000000000001100001010000
                ;mem[11858] <= 30'b000000000000000001100111110000
                ;mem[11859] <= 30'b000000000000000001101000000000
                ;mem[11860] <= 30'b000000000000000001101000010000
                ;mem[11861] <= 30'b000000000000000000110011010000
                ;mem[11862] <= 30'b000000000000000000110011100000
                ;mem[11863] <= 30'b000000000000000000110011110000
                ;mem[11864] <= 30'b000000000000000000110100000000
                ;mem[11865] <= 30'b000000000000000000110100010000
                ;mem[11866] <= 30'b000000000000000000111010000000
                ;mem[11867] <= 30'b000000000000000000111010010000
                ;mem[11868] <= 30'b000000000000000000111010100000
                ;mem[11869] <= 30'b000000000000000000111010110000
                ;mem[11870] <= 30'b000000000000000000111011000000
                ;mem[11871] <= 30'b000000000000000000111011010000
                ;mem[11872] <= 30'b000000000000000000111011100000
                ;mem[11873] <= 30'b000000000000000000111011110000
                ;mem[11874] <= 30'b000000000000000000111100000000
                ;mem[11875] <= 30'b000000000000000000111100010000
                ;mem[11876] <= 30'b000000000000000000111100100000
                ;mem[11877] <= 30'b000000000000000000111100110000
                ;mem[11878] <= 30'b000000001000000000000111010000
                ;mem[11879] <= 30'b000000001000000000000111100000
                ;mem[11880] <= 30'b000000001000000000000111110000
                ;mem[11881] <= 30'b000000001000000000001000000000
                ;mem[11882] <= 30'b000000001000000000001000010000
                ;mem[11883] <= 30'b000000001000000000001110000000
                ;mem[11884] <= 30'b000000001000000000001110010000
                ;mem[11885] <= 30'b000000001000000000001110100000
                ;mem[11886] <= 30'b000000001000000000001110110000
                ;mem[11887] <= 30'b000000001000000000001111000000
                ;mem[11888] <= 30'b000000001000000000001111010000
                ;mem[11889] <= 30'b000000001000000000001111100000
                ;mem[11890] <= 30'b000000001000000000001111110000
                ;mem[11891] <= 30'b000000001000000000010000000000
                ;mem[11892] <= 30'b000000001000000000010000010000
                ;mem[11893] <= 30'b000000001000000000010000100000
                ;mem[11894] <= 30'b000000001000000000010000110000
                ;mem[11895] <= 30'b000000001000000000010101000000
                ;mem[11896] <= 30'b000000001000000000010101010000
                ;mem[11897] <= 30'b000000001000000000010101100000
                ;mem[11898] <= 30'b000000001000000000010101110000
                ;mem[11899] <= 30'b000000001000000000010110000000
                ;mem[11900] <= 30'b000000001000000000010110010000
                ;mem[11901] <= 30'b000000001000000000010110100000
                ;mem[11902] <= 30'b000000001000000000010110110000
                ;mem[11903] <= 30'b000000001000000000010111000000
                ;mem[11904] <= 30'b000000001000000000010111010000
                ;mem[11905] <= 30'b000000001000000000010111100000
                ;mem[11906] <= 30'b000000001000000000010111110000
                ;mem[11907] <= 30'b000000001000000000011100010000
                ;mem[11908] <= 30'b000000001000000000011100100000
                ;mem[11909] <= 30'b000000001000000000011100110000
                ;mem[11910] <= 30'b000000001000000000011101000000
                ;mem[11911] <= 30'b000000001000000000011101010000
                ;mem[11912] <= 30'b000000001000000000011101100000
                ;mem[11913] <= 30'b000000001000000000011101110000
                ;mem[11914] <= 30'b000000001000000000011110000000
                ;mem[11915] <= 30'b000000001000000000011110010000
                ;mem[11916] <= 30'b000000001000000000011110100000
                ;mem[11917] <= 30'b000000001000000000011110110000
                ;mem[11918] <= 30'b000000001000000000100100110000
                ;mem[11919] <= 30'b000000001000000000100101000000
                ;mem[11920] <= 30'b000000001000000000100101010000
                ;mem[11921] <= 30'b000000001000000000100101100000
                ;mem[11922] <= 30'b000000001000000000100101110000
                ;mem[11923] <= 30'b000000001000000000101100000000
                ;mem[11924] <= 30'b000000001000000000101100010000
                ;mem[11925] <= 30'b000000001000000000101100100000
                ;mem[11926] <= 30'b000000001000000000101100110000
                ;mem[11927] <= 30'b000000001000000000110010110000
                ;mem[11928] <= 30'b000000001000000000110011000000
                ;mem[11929] <= 30'b000000001000000000110011010000
                ;mem[11930] <= 30'b000000001000000000110011100000
                ;mem[11931] <= 30'b000000001000000000111001100000
                ;mem[11932] <= 30'b000000001000000000111001110000
                ;mem[11933] <= 30'b000000001000000000111010000000
                ;mem[11934] <= 30'b000000001000000000111010010000
                ;mem[11935] <= 30'b000000001000000000111010100000
                ;mem[11936] <= 30'b000000010000000000000000000000
                ;mem[11937] <= 30'b000000010000000000000000010000
                ;mem[11938] <= 30'b000000010000000000000000100000
                ;mem[11939] <= 30'b000000010000000000000000110000
                ;mem[11940] <= 30'b000000010000000000000110110000
                ;mem[11941] <= 30'b000000010000000000000111000000
                ;mem[11942] <= 30'b000000010000000000000111010000
                ;mem[11943] <= 30'b000000010000000000000111100000
                ;mem[11944] <= 30'b000000010000000000001101100000
                ;mem[11945] <= 30'b000000010000000000001101110000
                ;mem[11946] <= 30'b000000010000000000001110000000
                ;mem[11947] <= 30'b000000010000000000001110010000
                ;mem[11948] <= 30'b000000010000000000001110100000
                ;mem[11949] <= 30'b000000010000000000010100100000
                ;mem[11950] <= 30'b000000010000000000010100110000
                ;mem[11951] <= 30'b000000010000000000010101000000
                ;mem[11952] <= 30'b000000010000000000010101010000
                ;mem[11953] <= 30'b000000010000000000011011010000
                ;mem[11954] <= 30'b000000010000000000011011100000
                ;mem[11955] <= 30'b000000010000000000011011110000
                ;mem[11956] <= 30'b000000010000000000011100000000
                ;mem[11957] <= 30'b000000010000000000100010010000
                ;mem[11958] <= 30'b000000010000000000100010100000
                ;mem[11959] <= 30'b000000010000000000100010110000
                ;mem[11960] <= 30'b000000010000000000100011000000
                ;mem[11961] <= 30'b000000010000000000101001000000
                ;mem[11962] <= 30'b000000010000000000101001010000
                ;mem[11963] <= 30'b000000010000000000101001100000
                ;mem[11964] <= 30'b000000010000000000101001110000
                ;mem[11965] <= 30'b000000010000000000101111110000
                ;mem[11966] <= 30'b000000010000000000110000000000
                ;mem[11967] <= 30'b000000010000000000110000010000
                ;mem[11968] <= 30'b000000010000000000110000100000
                ;mem[11969] <= 30'b000000010000000000110110110000
                ;mem[11970] <= 30'b000000010000000000110111000000
                ;mem[11971] <= 30'b000000010000000000110111010000
                ;mem[11972] <= 30'b000000010000000000110111100000
                ;mem[11973] <= 30'b000000010000000000111101110000
                ;mem[11974] <= 30'b000000010000000000111110000000
                ;mem[11975] <= 30'b000000010000000000111110010000
                ;mem[11976] <= 30'b000000010000000000111110100000
                ;mem[11977] <= 30'b000000000000000001000011110000
                ;mem[11978] <= 30'b000000000000000001000100000000
                ;mem[11979] <= 30'b000000000000000001000100010000
                ;mem[11980] <= 30'b000000000000000001000100100000
                ;mem[11981] <= 30'b000000000000000001001010110000
                ;mem[11982] <= 30'b000000000000000001001011000000
                ;mem[11983] <= 30'b000000000000000001001011010000
                ;mem[11984] <= 30'b000000000000000001001011100000
                ;mem[11985] <= 30'b000000000000000001010001110000
                ;mem[11986] <= 30'b000000000000000001010010000000
                ;mem[11987] <= 30'b000000000000000001010010010000
                ;mem[11988] <= 30'b000000000000000001010010100000
                ;mem[11989] <= 30'b000000000000000001011000110000
                ;mem[11990] <= 30'b000000000000000001011001000000
                ;mem[11991] <= 30'b000000000000000001011001010000
                ;mem[11992] <= 30'b000000000000000001011001100000
                ;mem[11993] <= 30'b000000000000000001011111110000
                ;mem[11994] <= 30'b000000000000000001100000000000
                ;mem[11995] <= 30'b000000000000000001100000010000
                ;mem[11996] <= 30'b000000000000000001100110100000
                ;mem[11997] <= 30'b000000000000000001100110110000
                ;mem[11998] <= 30'b000000000000000001100111000000
                ;mem[11999] <= 30'b000000000000000001100111010000
                ;mem[12000] <= 30'b000000000000000001101101110000
                ;mem[12001] <= 30'b000000000000000001101110000000
                ;mem[12002] <= 30'b000000000000000001110100110000
                ;mem[12003] <= 30'b000000000000000001110101000000
                ;mem[12004] <= 30'b000000000000000000100100110000
                ;mem[12005] <= 30'b000000000000000000100101000000
                ;mem[12006] <= 30'b000000000000000000100101010000
                ;mem[12007] <= 30'b000000000000000000100101100000
                ;mem[12008] <= 30'b000000000000000000100101110000
                ;mem[12009] <= 30'b000000000000000000100110000000
                ;mem[12010] <= 30'b000000000000000000100110010000
                ;mem[12011] <= 30'b000000000000000000100110100000
                ;mem[12012] <= 30'b000000000000000000101011100000
                ;mem[12013] <= 30'b000000000000000000101011110000
                ;mem[12014] <= 30'b000000000000000000101100000000
                ;mem[12015] <= 30'b000000000000000000101100010000
                ;mem[12016] <= 30'b000000000000000000101100100000
                ;mem[12017] <= 30'b000000000000000000101100110000
                ;mem[12018] <= 30'b000000000000000000101101000000
                ;mem[12019] <= 30'b000000000000000000101101010000
                ;mem[12020] <= 30'b000000000000000000101101100000
                ;mem[12021] <= 30'b000000000000000000110010010000
                ;mem[12022] <= 30'b000000000000000000110010100000
                ;mem[12023] <= 30'b000000000000000000110010110000
                ;mem[12024] <= 30'b000000000000000000110011000000
                ;mem[12025] <= 30'b000000000000000000110100010000
                ;mem[12026] <= 30'b000000000000000000110100100000
                ;mem[12027] <= 30'b000000000000000000111011010000
                ;mem[12028] <= 30'b000000000000000000111011100000
                ;mem[12029] <= 30'b000000001000000000000000000000
                ;mem[12030] <= 30'b000000001000000000000000010000
                ;mem[12031] <= 30'b000000001000000000000000100000
                ;mem[12032] <= 30'b000000001000000000000000110000
                ;mem[12033] <= 30'b000000001000000000000001000000
                ;mem[12034] <= 30'b000000001000000000000001010000
                ;mem[12035] <= 30'b000000001000000000000001100000
                ;mem[12036] <= 30'b000000001000000000000110010000
                ;mem[12037] <= 30'b000000001000000000000110100000
                ;mem[12038] <= 30'b000000001000000000000110110000
                ;mem[12039] <= 30'b000000001000000000000111000000
                ;mem[12040] <= 30'b000000001000000000001000010000
                ;mem[12041] <= 30'b000000001000000000001000100000
                ;mem[12042] <= 30'b000000001000000000001111010000
                ;mem[12043] <= 30'b000000001000000000001111100000
                ;mem[12044] <= 30'b000000001000000000010110000000
                ;mem[12045] <= 30'b000000001000000000010110010000
                ;mem[12046] <= 30'b000000001000000000010110100000
                ;mem[12047] <= 30'b000000001000000000011100110000
                ;mem[12048] <= 30'b000000001000000000011101000000
                ;mem[12049] <= 30'b000000001000000000011101010000
                ;mem[12050] <= 30'b000000001000000000100011100000
                ;mem[12051] <= 30'b000000001000000000100011110000
                ;mem[12052] <= 30'b000000001000000000100100000000
                ;mem[12053] <= 30'b000000001000000000100100010000
                ;mem[12054] <= 30'b000000001000000000101010010000
                ;mem[12055] <= 30'b000000001000000000101010100000
                ;mem[12056] <= 30'b000000001000000000101010110000
                ;mem[12057] <= 30'b000000001000000000101011000000
                ;mem[12058] <= 30'b000000001000000000101011010000
                ;mem[12059] <= 30'b000000001000000000101011100000
                ;mem[12060] <= 30'b000000001000000000101011110000
                ;mem[12061] <= 30'b000000001000000000101100000000
                ;mem[12062] <= 30'b000000001000000000110000110000
                ;mem[12063] <= 30'b000000001000000000110001000000
                ;mem[12064] <= 30'b000000001000000000110001010000
                ;mem[12065] <= 30'b000000001000000000110001100000
                ;mem[12066] <= 30'b000000001000000000110001110000
                ;mem[12067] <= 30'b000000001000000000110010010000
                ;mem[12068] <= 30'b000000001000000000110010100000
                ;mem[12069] <= 30'b000000001000000000110010110000
                ;mem[12070] <= 30'b000000001000000000110011000000
                ;mem[12071] <= 30'b000000001000000000110011010000
                ;mem[12072] <= 30'b000000001000000000111000000000
                ;mem[12073] <= 30'b000000001000000000111000010000
                ;mem[12074] <= 30'b000000001000000000111010000000
                ;mem[12075] <= 30'b000000001000000000111010010000
                ;mem[12076] <= 30'b000000001000000000111010100000
                ;mem[12077] <= 30'b000000001000000000111011110000
                ;mem[12078] <= 30'b000000010000000000000000000000
                ;mem[12079] <= 30'b000000010000000000000100110000
                ;mem[12080] <= 30'b000000010000000000000101000000
                ;mem[12081] <= 30'b000000010000000000000101010000
                ;mem[12082] <= 30'b000000010000000000000101100000
                ;mem[12083] <= 30'b000000010000000000000101110000
                ;mem[12084] <= 30'b000000010000000000000110010000
                ;mem[12085] <= 30'b000000010000000000000110100000
                ;mem[12086] <= 30'b000000010000000000000110110000
                ;mem[12087] <= 30'b000000010000000000000111000000
                ;mem[12088] <= 30'b000000010000000000000111010000
                ;mem[12089] <= 30'b000000010000000000001100000000
                ;mem[12090] <= 30'b000000010000000000001100010000
                ;mem[12091] <= 30'b000000010000000000001110000000
                ;mem[12092] <= 30'b000000010000000000001110010000
                ;mem[12093] <= 30'b000000010000000000001110100000
                ;mem[12094] <= 30'b000000010000000000001111110000
                ;mem[12095] <= 30'b000000010000000000010101010000
                ;mem[12096] <= 30'b000000010000000000010101100000
                ;mem[12097] <= 30'b000000010000000000010110010000
                ;mem[12098] <= 30'b000000010000000000010110100000
                ;mem[12099] <= 30'b000000010000000000011100100000
                ;mem[12100] <= 30'b000000010000000000011100110000
                ;mem[12101] <= 30'b000000010000000000011101000000
                ;mem[12102] <= 30'b000000010000000000011101010000
                ;mem[12103] <= 30'b000000010000000000100011100000
                ;mem[12104] <= 30'b000000010000000000100011110000
                ;mem[12105] <= 30'b000000010000000000100100000000
                ;mem[12106] <= 30'b000000010000000000101010000000
                ;mem[12107] <= 30'b000000010000000000101010010000
                ;mem[12108] <= 30'b000000010000000000101010100000
                ;mem[12109] <= 30'b000000010000000000101010110000
                ;mem[12110] <= 30'b000000010000000000110000110000
                ;mem[12111] <= 30'b000000010000000000110001000000
                ;mem[12112] <= 30'b000000010000000000110001010000
                ;mem[12113] <= 30'b000000010000000000110001100000
                ;mem[12114] <= 30'b000000010000000000110001110000
                ;mem[12115] <= 30'b000000010000000000110111100000
                ;mem[12116] <= 30'b000000010000000000110111110000
                ;mem[12117] <= 30'b000000010000000000111000010000
                ;mem[12118] <= 30'b000000010000000000111000100000
                ;mem[12119] <= 30'b000000010000000000111000110000
                ;mem[12120] <= 30'b000000010000000000111110010000
                ;mem[12121] <= 30'b000000010000000000111110100000
                ;mem[12122] <= 30'b000000010000000000111111000000
                ;mem[12123] <= 30'b000000010000000000111111010000
                ;mem[12124] <= 30'b000000010000000000111111100000
                ;mem[12125] <= 30'b000000000000000001000100110000
                ;mem[12126] <= 30'b000000000000000001000101000000
                ;mem[12127] <= 30'b000000000000000001000101010000
                ;mem[12128] <= 30'b000000000000000001000101100000
                ;mem[12129] <= 30'b000000000000000001000101110000
                ;mem[12130] <= 30'b000000000000000001001011100000
                ;mem[12131] <= 30'b000000000000000001001011110000
                ;mem[12132] <= 30'b000000000000000001001100010000
                ;mem[12133] <= 30'b000000000000000001001100100000
                ;mem[12134] <= 30'b000000000000000001001100110000
                ;mem[12135] <= 30'b000000000000000001010010010000
                ;mem[12136] <= 30'b000000000000000001010010100000
                ;mem[12137] <= 30'b000000000000000001010011000000
                ;mem[12138] <= 30'b000000000000000001010011010000
                ;mem[12139] <= 30'b000000000000000001010011100000
                ;mem[12140] <= 30'b000000000000000001011001000000
                ;mem[12141] <= 30'b000000000000000001011001010000
                ;mem[12142] <= 30'b000000000000000001011001110000
                ;mem[12143] <= 30'b000000000000000001011010000000
                ;mem[12144] <= 30'b000000000000000001011010010000
                ;mem[12145] <= 30'b000000000000000001011010100000
                ;mem[12146] <= 30'b000000000000000001100000000000
                ;mem[12147] <= 30'b000000000000000001100000010000
                ;mem[12148] <= 30'b000000000000000001100000100000
                ;mem[12149] <= 30'b000000000000000001100000110000
                ;mem[12150] <= 30'b000000000000000001100001000000
                ;mem[12151] <= 30'b000000000000000001100001010000
                ;mem[12152] <= 30'b000000000000000001100111000000
                ;mem[12153] <= 30'b000000000000000001100111010000
                ;mem[12154] <= 30'b000000000000000001100111100000
                ;mem[12155] <= 30'b000000000000000001100111110000
                ;mem[12156] <= 30'b000000000000000000010001000000
                ;mem[12157] <= 30'b000000000000000000010001010000
                ;mem[12158] <= 30'b000000000000000000010111110000
                ;mem[12159] <= 30'b000000000000000000011000000000
                ;mem[12160] <= 30'b000000000000000000011000010000
                ;mem[12161] <= 30'b000000000000000000011000100000
                ;mem[12162] <= 30'b000000000000000000011110110000
                ;mem[12163] <= 30'b000000000000000000011111000000
                ;mem[12164] <= 30'b000000000000000000011111100000
                ;mem[12165] <= 30'b000000000000000000100101100000
                ;mem[12166] <= 30'b000000000000000000100101110000
                ;mem[12167] <= 30'b000000000000000000100110000000
                ;mem[12168] <= 30'b000000000000000000101100100000
                ;mem[12169] <= 30'b000000000000000000101100110000
                ;mem[12170] <= 30'b000000000000000000110011010000
                ;mem[12171] <= 30'b000000000000000000110011100000
                ;mem[12172] <= 30'b000000000000000000110011110000
                ;mem[12173] <= 30'b000000000000000000111010010000
                ;mem[12174] <= 30'b000000000000000000111010100000
                ;mem[12175] <= 30'b000000001000000000000000100000
                ;mem[12176] <= 30'b000000001000000000000000110000
                ;mem[12177] <= 30'b000000001000000000000111010000
                ;mem[12178] <= 30'b000000001000000000000111100000
                ;mem[12179] <= 30'b000000001000000000000111110000
                ;mem[12180] <= 30'b000000001000000000001110010000
                ;mem[12181] <= 30'b000000001000000000001110100000
                ;mem[12182] <= 30'b000000001000000000010101010000
                ;mem[12183] <= 30'b000000001000000000010101100000
                ;mem[12184] <= 30'b000000001000000000011100000000
                ;mem[12185] <= 30'b000000001000000000011100010000
                ;mem[12186] <= 30'b000000001000000000011100100000
                ;mem[12187] <= 30'b000000001000000000100011000000
                ;mem[12188] <= 30'b000000001000000000100011010000
                ;mem[12189] <= 30'b000000001000000000100011100000
                ;mem[12190] <= 30'b000000001000000000100101110000
                ;mem[12191] <= 30'b000000001000000000100110000000
                ;mem[12192] <= 30'b000000001000000000101010000000
                ;mem[12193] <= 30'b000000001000000000101010010000
                ;mem[12194] <= 30'b000000001000000000101010100000
                ;mem[12195] <= 30'b000000001000000000101100100000
                ;mem[12196] <= 30'b000000001000000000101100110000
                ;mem[12197] <= 30'b000000001000000000101101000000
                ;mem[12198] <= 30'b000000001000000000101101010000
                ;mem[12199] <= 30'b000000001000000000110001000000
                ;mem[12200] <= 30'b000000001000000000110001010000
                ;mem[12201] <= 30'b000000001000000000110001100000
                ;mem[12202] <= 30'b000000001000000000110011010000
                ;mem[12203] <= 30'b000000001000000000110011100000
                ;mem[12204] <= 30'b000000001000000000110011110000
                ;mem[12205] <= 30'b000000001000000000110100000000
                ;mem[12206] <= 30'b000000001000000000110100010000
                ;mem[12207] <= 30'b000000001000000000110100100000
                ;mem[12208] <= 30'b000000001000000000111000000000
                ;mem[12209] <= 30'b000000001000000000111000010000
                ;mem[12210] <= 30'b000000001000000000111000100000
                ;mem[12211] <= 30'b000000001000000000111010000000
                ;mem[12212] <= 30'b000000001000000000111010010000
                ;mem[12213] <= 30'b000000001000000000111010100000
                ;mem[12214] <= 30'b000000001000000000111010110000
                ;mem[12215] <= 30'b000000001000000000111011010000
                ;mem[12216] <= 30'b000000001000000000111011100000
                ;mem[12217] <= 30'b000000001000000000111111010000
                ;mem[12218] <= 30'b000000001000000000111111100000
                ;mem[12219] <= 30'b000000010000000000000000100000
                ;mem[12220] <= 30'b000000010000000000000000110000
                ;mem[12221] <= 30'b000000010000000000000001000000
                ;mem[12222] <= 30'b000000010000000000000001010000
                ;mem[12223] <= 30'b000000010000000000000101000000
                ;mem[12224] <= 30'b000000010000000000000101010000
                ;mem[12225] <= 30'b000000010000000000000101100000
                ;mem[12226] <= 30'b000000010000000000000111010000
                ;mem[12227] <= 30'b000000010000000000000111100000
                ;mem[12228] <= 30'b000000010000000000000111110000
                ;mem[12229] <= 30'b000000010000000000001000000000
                ;mem[12230] <= 30'b000000010000000000001000010000
                ;mem[12231] <= 30'b000000010000000000001000100000
                ;mem[12232] <= 30'b000000010000000000001100000000
                ;mem[12233] <= 30'b000000010000000000001100010000
                ;mem[12234] <= 30'b000000010000000000001100100000
                ;mem[12235] <= 30'b000000010000000000001110000000
                ;mem[12236] <= 30'b000000010000000000001110010000
                ;mem[12237] <= 30'b000000010000000000001110100000
                ;mem[12238] <= 30'b000000010000000000001110110000
                ;mem[12239] <= 30'b000000010000000000001111010000
                ;mem[12240] <= 30'b000000010000000000001111100000
                ;mem[12241] <= 30'b000000010000000000010011010000
                ;mem[12242] <= 30'b000000010000000000010011100000
                ;mem[12243] <= 30'b000000010000000000010100110000
                ;mem[12244] <= 30'b000000010000000000010101000000
                ;mem[12245] <= 30'b000000010000000000010101010000
                ;mem[12246] <= 30'b000000010000000000010110010000
                ;mem[12247] <= 30'b000000010000000000010110100000
                ;mem[12248] <= 30'b000000010000000000010110110000
                ;mem[12249] <= 30'b000000010000000000011010010000
                ;mem[12250] <= 30'b000000010000000000011010100000
                ;mem[12251] <= 30'b000000010000000000011011100000
                ;mem[12252] <= 30'b000000010000000000011011110000
                ;mem[12253] <= 30'b000000010000000000011100000000
                ;mem[12254] <= 30'b000000010000000000011101010000
                ;mem[12255] <= 30'b000000010000000000011101100000
                ;mem[12256] <= 30'b000000010000000000011101110000
                ;mem[12257] <= 30'b000000010000000000100001010000
                ;mem[12258] <= 30'b000000010000000000100001100000
                ;mem[12259] <= 30'b000000010000000000100001110000
                ;mem[12260] <= 30'b000000010000000000100010100000
                ;mem[12261] <= 30'b000000010000000000100010110000
                ;mem[12262] <= 30'b000000010000000000100100010000
                ;mem[12263] <= 30'b000000010000000000100100100000
                ;mem[12264] <= 30'b000000010000000000101000100000
                ;mem[12265] <= 30'b000000010000000000101000110000
                ;mem[12266] <= 30'b000000010000000000101001000000
                ;mem[12267] <= 30'b000000010000000000101001010000
                ;mem[12268] <= 30'b000000010000000000101001100000
                ;mem[12269] <= 30'b000000010000000000101001110000
                ;mem[12270] <= 30'b000000010000000000101010110000
                ;mem[12271] <= 30'b000000010000000000101011000000
                ;mem[12272] <= 30'b000000010000000000101011010000
                ;mem[12273] <= 30'b000000010000000000101011100000
                ;mem[12274] <= 30'b000000010000000000101111110000
                ;mem[12275] <= 30'b000000010000000000110000000000
                ;mem[12276] <= 30'b000000010000000000110000010000
                ;mem[12277] <= 30'b000000010000000000110000100000
                ;mem[12278] <= 30'b000000010000000000110000110000
                ;mem[12279] <= 30'b000000010000000000110001000000
                ;mem[12280] <= 30'b000000010000000000110001010000
                ;mem[12281] <= 30'b000000010000000000110001100000
                ;mem[12282] <= 30'b000000010000000000110001110000
                ;mem[12283] <= 30'b000000010000000000110010000000
                ;mem[12284] <= 30'b000000010000000000110010010000
                ;mem[12285] <= 30'b000000010000000000110111000000
                ;mem[12286] <= 30'b000000010000000000110111010000
                ;mem[12287] <= 30'b000000010000000000110111100000
                ;mem[12288] <= 30'b000000010000000000110111110000
                ;mem[12289] <= 30'b000000010000000000111000000000
                ;mem[12290] <= 30'b000000010000000000111000010000
                ;mem[12291] <= 30'b000000010000000000111000100000
                ;mem[12292] <= 30'b000000010000000000111000110000
                ;mem[12293] <= 30'b000000010000000000111110100000
                ;mem[12294] <= 30'b000000010000000000111110110000
                ;mem[12295] <= 30'b000000010000000000111111000000
                ;mem[12296] <= 30'b000000010000000000111111010000
                ;mem[12297] <= 30'b000000010000000000111111100000
                ;mem[12298] <= 30'b000000000000000001000011110000
                ;mem[12299] <= 30'b000000000000000001000100000000
                ;mem[12300] <= 30'b000000000000000001000100010000
                ;mem[12301] <= 30'b000000000000000001000100100000
                ;mem[12302] <= 30'b000000000000000001000100110000
                ;mem[12303] <= 30'b000000000000000001000101000000
                ;mem[12304] <= 30'b000000000000000001000101010000
                ;mem[12305] <= 30'b000000000000000001000101100000
                ;mem[12306] <= 30'b000000000000000001000101110000
                ;mem[12307] <= 30'b000000000000000001000110000000
                ;mem[12308] <= 30'b000000000000000001000110010000
                ;mem[12309] <= 30'b000000000000000001001011000000
                ;mem[12310] <= 30'b000000000000000001001011010000
                ;mem[12311] <= 30'b000000000000000001001011100000
                ;mem[12312] <= 30'b000000000000000001001011110000
                ;mem[12313] <= 30'b000000000000000001001100000000
                ;mem[12314] <= 30'b000000000000000001001100010000
                ;mem[12315] <= 30'b000000000000000001001100100000
                ;mem[12316] <= 30'b000000000000000001001100110000
                ;mem[12317] <= 30'b000000000000000001010010100000
                ;mem[12318] <= 30'b000000000000000001010010110000
                ;mem[12319] <= 30'b000000000000000001010011000000
                ;mem[12320] <= 30'b000000000000000001010011010000
                ;mem[12321] <= 30'b000000000000000001010011100000
                ;mem[12322] <= 30'b000000000000000000100000010000
                ;mem[12323] <= 30'b000000000000000000100000100000
                ;mem[12324] <= 30'b000000000000000000100111010000
                ;mem[12325] <= 30'b000000000000000000100111100000
                ;mem[12326] <= 30'b000000000000000000101110010000
                ;mem[12327] <= 30'b000000000000000000101110100000
                ;mem[12328] <= 30'b000000000000000000110101000000
                ;mem[12329] <= 30'b000000000000000000110101010000
                ;mem[12330] <= 30'b000000000000000000110101100000
                ;mem[12331] <= 30'b000000000000000000111011110000
                ;mem[12332] <= 30'b000000000000000000111100000000
                ;mem[12333] <= 30'b000000000000000000111100010000
                ;mem[12334] <= 30'b000000000000000000111100100000
                ;mem[12335] <= 30'b000000001000000000000010010000
                ;mem[12336] <= 30'b000000001000000000000010100000
                ;mem[12337] <= 30'b000000001000000000001001000000
                ;mem[12338] <= 30'b000000001000000000001001010000
                ;mem[12339] <= 30'b000000001000000000001001100000
                ;mem[12340] <= 30'b000000001000000000001111110000
                ;mem[12341] <= 30'b000000001000000000010000000000
                ;mem[12342] <= 30'b000000001000000000010000010000
                ;mem[12343] <= 30'b000000001000000000010000100000
                ;mem[12344] <= 30'b000000001000000000010110110000
                ;mem[12345] <= 30'b000000001000000000010111000000
                ;mem[12346] <= 30'b000000001000000000010111010000
                ;mem[12347] <= 30'b000000001000000000011101100000
                ;mem[12348] <= 30'b000000001000000000011101110000
                ;mem[12349] <= 30'b000000001000000000011110000000
                ;mem[12350] <= 30'b000000001000000000100100100000
                ;mem[12351] <= 30'b000000001000000000100100110000
                ;mem[12352] <= 30'b000000001000000000100101000000
                ;mem[12353] <= 30'b000000001000000000101011010000
                ;mem[12354] <= 30'b000000001000000000101011100000
                ;mem[12355] <= 30'b000000001000000000101011110000
                ;mem[12356] <= 30'b000000001000000000101100000000
                ;mem[12357] <= 30'b000000001000000000110010010000
                ;mem[12358] <= 30'b000000001000000000110010100000
                ;mem[12359] <= 30'b000000001000000000110010110000
                ;mem[12360] <= 30'b000000001000000000110011000000
                ;mem[12361] <= 30'b000000001000000000111001000000
                ;mem[12362] <= 30'b000000001000000000111001010000
                ;mem[12363] <= 30'b000000001000000000111001100000
                ;mem[12364] <= 30'b000000001000000000111001110000
                ;mem[12365] <= 30'b000000010000000000000000000000
                ;mem[12366] <= 30'b000000010000000000000110010000
                ;mem[12367] <= 30'b000000010000000000000110100000
                ;mem[12368] <= 30'b000000010000000000000110110000
                ;mem[12369] <= 30'b000000010000000000000111000000
                ;mem[12370] <= 30'b000000010000000000001101000000
                ;mem[12371] <= 30'b000000010000000000001101010000
                ;mem[12372] <= 30'b000000010000000000001101100000
                ;mem[12373] <= 30'b000000010000000000001101110000
                ;mem[12374] <= 30'b000000010000000000010100000000
                ;mem[12375] <= 30'b000000010000000000010100010000
                ;mem[12376] <= 30'b000000010000000000010100100000
                ;mem[12377] <= 30'b000000010000000000010100110000
                ;mem[12378] <= 30'b000000010000000000011011010000
                ;mem[12379] <= 30'b000000010000000000011011100000
                ;mem[12380] <= 30'b000000010000000000011011110000
                ;mem[12381] <= 30'b000000010000000000011100000000
                ;mem[12382] <= 30'b000000010000000000100010000000
                ;mem[12383] <= 30'b000000010000000000100010010000
                ;mem[12384] <= 30'b000000010000000000100010100000
                ;mem[12385] <= 30'b000000010000000000100010110000
                ;mem[12386] <= 30'b000000010000000000101001000000
                ;mem[12387] <= 30'b000000010000000000101001010000
                ;mem[12388] <= 30'b000000010000000000101001100000
                ;mem[12389] <= 30'b000000010000000000101111110000
                ;mem[12390] <= 30'b000000010000000000110000000000
                ;mem[12391] <= 30'b000000010000000000110000010000
                ;mem[12392] <= 30'b000000010000000000110000100000
                ;mem[12393] <= 30'b000000010000000000110110100000
                ;mem[12394] <= 30'b000000010000000000110110110000
                ;mem[12395] <= 30'b000000010000000000110111000000
                ;mem[12396] <= 30'b000000010000000000110111010000
                ;mem[12397] <= 30'b000000010000000000110111100000
                ;mem[12398] <= 30'b000000010000000000111101100000
                ;mem[12399] <= 30'b000000010000000000111101110000
                ;mem[12400] <= 30'b000000010000000000111110000000
                ;mem[12401] <= 30'b000000010000000000111110010000
                ;mem[12402] <= 30'b000000000000000001000011110000
                ;mem[12403] <= 30'b000000000000000001000100000000
                ;mem[12404] <= 30'b000000000000000001000100010000
                ;mem[12405] <= 30'b000000000000000001000100100000
                ;mem[12406] <= 30'b000000000000000001001010100000
                ;mem[12407] <= 30'b000000000000000001001010110000
                ;mem[12408] <= 30'b000000000000000001001011000000
                ;mem[12409] <= 30'b000000000000000001001011010000
                ;mem[12410] <= 30'b000000000000000001001011100000
                ;mem[12411] <= 30'b000000000000000001010001100000
                ;mem[12412] <= 30'b000000000000000001010001110000
                ;mem[12413] <= 30'b000000000000000001010010000000
                ;mem[12414] <= 30'b000000000000000001010010010000
                ;mem[12415] <= 30'b000000000000000001011000100000
                ;mem[12416] <= 30'b000000000000000001011000110000
                ;mem[12417] <= 30'b000000000000000001011001000000
                ;mem[12418] <= 30'b000000000000000001011001010000
                ;mem[12419] <= 30'b000000000000000001100000000000
                ;mem[12420] <= 30'b000000000000000000100110100000
                ;mem[12421] <= 30'b000000000000000000100110110000
                ;mem[12422] <= 30'b000000000000000000100111000000
                ;mem[12423] <= 30'b000000000000000000100111010000
                ;mem[12424] <= 30'b000000000000000000100111100000
                ;mem[12425] <= 30'b000000000000000000101101000000
                ;mem[12426] <= 30'b000000000000000000101101010000
                ;mem[12427] <= 30'b000000000000000000101101100000
                ;mem[12428] <= 30'b000000000000000000101101110000
                ;mem[12429] <= 30'b000000000000000000101110000000
                ;mem[12430] <= 30'b000000000000000000101110010000
                ;mem[12431] <= 30'b000000000000000000101110100000
                ;mem[12432] <= 30'b000000000000000000101110110000
                ;mem[12433] <= 30'b000000000000000000110011100000
                ;mem[12434] <= 30'b000000000000000000110011110000
                ;mem[12435] <= 30'b000000000000000000110100000000
                ;mem[12436] <= 30'b000000000000000000110100010000
                ;mem[12437] <= 30'b000000000000000000110100100000
                ;mem[12438] <= 30'b000000000000000000110101100000
                ;mem[12439] <= 30'b000000000000000000110101110000
                ;mem[12440] <= 30'b000000000000000000111010100000
                ;mem[12441] <= 30'b000000000000000000111010110000
                ;mem[12442] <= 30'b000000000000000000111011000000
                ;mem[12443] <= 30'b000000000000000000111100100000
                ;mem[12444] <= 30'b000000000000000000111100110000
                ;mem[12445] <= 30'b000000001000000000000001000000
                ;mem[12446] <= 30'b000000001000000000000001010000
                ;mem[12447] <= 30'b000000001000000000000001100000
                ;mem[12448] <= 30'b000000001000000000000001110000
                ;mem[12449] <= 30'b000000001000000000000010000000
                ;mem[12450] <= 30'b000000001000000000000010010000
                ;mem[12451] <= 30'b000000001000000000000010100000
                ;mem[12452] <= 30'b000000001000000000000010110000
                ;mem[12453] <= 30'b000000001000000000000111100000
                ;mem[12454] <= 30'b000000001000000000000111110000
                ;mem[12455] <= 30'b000000001000000000001000000000
                ;mem[12456] <= 30'b000000001000000000001000010000
                ;mem[12457] <= 30'b000000001000000000001000100000
                ;mem[12458] <= 30'b000000001000000000001001100000
                ;mem[12459] <= 30'b000000001000000000001001110000
                ;mem[12460] <= 30'b000000001000000000001110100000
                ;mem[12461] <= 30'b000000001000000000001110110000
                ;mem[12462] <= 30'b000000001000000000001111000000
                ;mem[12463] <= 30'b000000001000000000010000100000
                ;mem[12464] <= 30'b000000001000000000010000110000
                ;mem[12465] <= 30'b000000001000000000010101100000
                ;mem[12466] <= 30'b000000001000000000010111010000
                ;mem[12467] <= 30'b000000001000000000010111100000
                ;mem[12468] <= 30'b000000001000000000011101110000
                ;mem[12469] <= 30'b000000001000000000011110000000
                ;mem[12470] <= 30'b000000001000000000011110010000
                ;mem[12471] <= 30'b000000001000000000011110100000
                ;mem[12472] <= 30'b000000001000000000100100100000
                ;mem[12473] <= 30'b000000001000000000100100110000
                ;mem[12474] <= 30'b000000001000000000100101000000
                ;mem[12475] <= 30'b000000001000000000100101010000
                ;mem[12476] <= 30'b000000001000000000101010110000
                ;mem[12477] <= 30'b000000001000000000101011000000
                ;mem[12478] <= 30'b000000001000000000101011010000
                ;mem[12479] <= 30'b000000001000000000101011100000
                ;mem[12480] <= 30'b000000001000000000101011110000
                ;mem[12481] <= 30'b000000001000000000101100000000
                ;mem[12482] <= 30'b000000001000000000101100010000
                ;mem[12483] <= 30'b000000001000000000110001110000
                ;mem[12484] <= 30'b000000001000000000110010000000
                ;mem[12485] <= 30'b000000001000000000110010010000
                ;mem[12486] <= 30'b000000001000000000110010100000
                ;mem[12487] <= 30'b000000001000000000110010110000
                ;mem[12488] <= 30'b000000001000000000110011000000
                ;mem[12489] <= 30'b000000001000000000110011010000
                ;mem[12490] <= 30'b000000001000000000110011100000
                ;mem[12491] <= 30'b000000001000000000111010010000
                ;mem[12492] <= 30'b000000001000000000111010100000
                ;mem[12493] <= 30'b000000001000000000111010110000
                ;mem[12494] <= 30'b000000010000000000000000000000
                ;mem[12495] <= 30'b000000010000000000000000010000
                ;mem[12496] <= 30'b000000010000000000000101110000
                ;mem[12497] <= 30'b000000010000000000000110000000
                ;mem[12498] <= 30'b000000010000000000000110010000
                ;mem[12499] <= 30'b000000010000000000000110100000
                ;mem[12500] <= 30'b000000010000000000000110110000
                ;mem[12501] <= 30'b000000010000000000000111000000
                ;mem[12502] <= 30'b000000010000000000000111010000
                ;mem[12503] <= 30'b000000010000000000000111100000
                ;mem[12504] <= 30'b000000010000000000001110010000
                ;mem[12505] <= 30'b000000010000000000001110100000
                ;mem[12506] <= 30'b000000010000000000001110110000
                ;mem[12507] <= 30'b000000010000000000010101100000
                ;mem[12508] <= 30'b000000010000000000010101110000
                ;mem[12509] <= 30'b000000010000000000011100110000
                ;mem[12510] <= 30'b000000010000000000011101000000
                ;mem[12511] <= 30'b000000010000000000100011100000
                ;mem[12512] <= 30'b000000010000000000100011110000
                ;mem[12513] <= 30'b000000010000000000100100000000
                ;mem[12514] <= 30'b000000010000000000101010100000
                ;mem[12515] <= 30'b000000010000000000101010110000
                ;mem[12516] <= 30'b000000010000000000101110110000
                ;mem[12517] <= 30'b000000010000000000101111000000
                ;mem[12518] <= 30'b000000010000000000110001100000
                ;mem[12519] <= 30'b000000010000000000110001110000
                ;mem[12520] <= 30'b000000010000000000110101110000
                ;mem[12521] <= 30'b000000010000000000110110000000
                ;mem[12522] <= 30'b000000010000000000111000010000
                ;mem[12523] <= 30'b000000010000000000111000100000
                ;mem[12524] <= 30'b000000010000000000111000110000
                ;mem[12525] <= 30'b000000010000000000111100110000
                ;mem[12526] <= 30'b000000010000000000111101000000
                ;mem[12527] <= 30'b000000010000000000111110110000
                ;mem[12528] <= 30'b000000010000000000111111000000
                ;mem[12529] <= 30'b000000010000000000111111010000
                ;mem[12530] <= 30'b000000010000000000111111100000
                ;mem[12531] <= 30'b000000000000000001000010110000
                ;mem[12532] <= 30'b000000000000000001000011000000
                ;mem[12533] <= 30'b000000000000000001000101100000
                ;mem[12534] <= 30'b000000000000000001000101110000
                ;mem[12535] <= 30'b000000000000000001001001110000
                ;mem[12536] <= 30'b000000000000000001001010000000
                ;mem[12537] <= 30'b000000000000000001001100010000
                ;mem[12538] <= 30'b000000000000000001001100100000
                ;mem[12539] <= 30'b000000000000000001001100110000
                ;mem[12540] <= 30'b000000000000000001010000110000
                ;mem[12541] <= 30'b000000000000000001010001000000
                ;mem[12542] <= 30'b000000000000000001010010110000
                ;mem[12543] <= 30'b000000000000000001010011000000
                ;mem[12544] <= 30'b000000000000000001010011010000
                ;mem[12545] <= 30'b000000000000000001010011100000
                ;mem[12546] <= 30'b000000000000000001010111110000
                ;mem[12547] <= 30'b000000000000000001011000000000
                ;mem[12548] <= 30'b000000000000000001011000010000
                ;mem[12549] <= 30'b000000000000000001011001010000
                ;mem[12550] <= 30'b000000000000000001011001100000
                ;mem[12551] <= 30'b000000000000000001011001110000
                ;mem[12552] <= 30'b000000000000000001011010000000
                ;mem[12553] <= 30'b000000000000000001011010010000
                ;mem[12554] <= 30'b000000000000000001011110110000
                ;mem[12555] <= 30'b000000000000000001011111000000
                ;mem[12556] <= 30'b000000000000000001011111010000
                ;mem[12557] <= 30'b000000000000000001011111100000
                ;mem[12558] <= 30'b000000000000000001011111110000
                ;mem[12559] <= 30'b000000000000000001100000000000
                ;mem[12560] <= 30'b000000000000000001100000010000
                ;mem[12561] <= 30'b000000000000000001100000100000
                ;mem[12562] <= 30'b000000000000000001100000110000
                ;mem[12563] <= 30'b000000000000000001100110010000
                ;mem[12564] <= 30'b000000000000000001100110100000
                ;mem[12565] <= 30'b000000000000000001100110110000
                ;mem[12566] <= 30'b000000000000000001100111000000
                ;mem[12567] <= 30'b000000000000000001100111010000
                ;mem[12568] <= 30'b000000000000000000010010000000
                ;mem[12569] <= 30'b000000000000000000010010010000
                ;mem[12570] <= 30'b000000000000000000011000110000
                ;mem[12571] <= 30'b000000000000000000011001000000
                ;mem[12572] <= 30'b000000000000000000011001010000
                ;mem[12573] <= 30'b000000000000000000011111110000
                ;mem[12574] <= 30'b000000000000000000100000000000
                ;mem[12575] <= 30'b000000000000000000100110100000
                ;mem[12576] <= 30'b000000000000000000100110110000
                ;mem[12577] <= 30'b000000000000000000101101010000
                ;mem[12578] <= 30'b000000000000000000101101100000
                ;mem[12579] <= 30'b000000000000000000110100010000
                ;mem[12580] <= 30'b000000000000000000110100100000
                ;mem[12581] <= 30'b000000000000000000111011000000
                ;mem[12582] <= 30'b000000000000000000111011010000
                ;mem[12583] <= 30'b000000001000000000000001010000
                ;mem[12584] <= 30'b000000001000000000000001100000
                ;mem[12585] <= 30'b000000001000000000001000010000
                ;mem[12586] <= 30'b000000001000000000001000100000
                ;mem[12587] <= 30'b000000001000000000001111000000
                ;mem[12588] <= 30'b000000001000000000001111010000
                ;mem[12589] <= 30'b000000001000000000010101110000
                ;mem[12590] <= 30'b000000001000000000010110000000
                ;mem[12591] <= 30'b000000001000000000011100100000
                ;mem[12592] <= 30'b000000001000000000011100110000
                ;mem[12593] <= 30'b000000001000000000011101000000
                ;mem[12594] <= 30'b000000001000000000100011100000
                ;mem[12595] <= 30'b000000001000000000100011110000
                ;mem[12596] <= 30'b000000001000000000101010100000
                ;mem[12597] <= 30'b000000001000000000101010110000
                ;mem[12598] <= 30'b000000001000000000110001010000
                ;mem[12599] <= 30'b000000001000000000110001100000
                ;mem[12600] <= 30'b000000001000000000110001110000
                ;mem[12601] <= 30'b000000001000000000110010110000
                ;mem[12602] <= 30'b000000001000000000110011000000
                ;mem[12603] <= 30'b000000001000000000110011010000
                ;mem[12604] <= 30'b000000001000000000110011100000
                ;mem[12605] <= 30'b000000001000000000110011110000
                ;mem[12606] <= 30'b000000001000000000111000010000
                ;mem[12607] <= 30'b000000001000000000111000100000
                ;mem[12608] <= 30'b000000001000000000111000110000
                ;mem[12609] <= 30'b000000001000000000111001100000
                ;mem[12610] <= 30'b000000001000000000111001110000
                ;mem[12611] <= 30'b000000001000000000111010000000
                ;mem[12612] <= 30'b000000001000000000111010100000
                ;mem[12613] <= 30'b000000001000000000111010110000
                ;mem[12614] <= 30'b000000001000000000111111010000
                ;mem[12615] <= 30'b000000001000000000111111100000
                ;mem[12616] <= 30'b000000001000000000111111110000
                ;mem[12617] <= 30'b000000010000000000000101010000
                ;mem[12618] <= 30'b000000010000000000000101100000
                ;mem[12619] <= 30'b000000010000000000000101110000
                ;mem[12620] <= 30'b000000010000000000000110110000
                ;mem[12621] <= 30'b000000010000000000000111000000
                ;mem[12622] <= 30'b000000010000000000000111010000
                ;mem[12623] <= 30'b000000010000000000000111100000
                ;mem[12624] <= 30'b000000010000000000000111110000
                ;mem[12625] <= 30'b000000010000000000001100010000
                ;mem[12626] <= 30'b000000010000000000001100100000
                ;mem[12627] <= 30'b000000010000000000001100110000
                ;mem[12628] <= 30'b000000010000000000001101100000
                ;mem[12629] <= 30'b000000010000000000001101110000
                ;mem[12630] <= 30'b000000010000000000001110000000
                ;mem[12631] <= 30'b000000010000000000001110100000
                ;mem[12632] <= 30'b000000010000000000001110110000
                ;mem[12633] <= 30'b000000010000000000010011010000
                ;mem[12634] <= 30'b000000010000000000010011100000
                ;mem[12635] <= 30'b000000010000000000010011110000
                ;mem[12636] <= 30'b000000010000000000010100010000
                ;mem[12637] <= 30'b000000010000000000010100100000
                ;mem[12638] <= 30'b000000010000000000010100110000
                ;mem[12639] <= 30'b000000010000000000010101100000
                ;mem[12640] <= 30'b000000010000000000010101110000
                ;mem[12641] <= 30'b000000010000000000010110000000
                ;mem[12642] <= 30'b000000010000000000011010010000
                ;mem[12643] <= 30'b000000010000000000011010100000
                ;mem[12644] <= 30'b000000010000000000011010110000
                ;mem[12645] <= 30'b000000010000000000011011000000
                ;mem[12646] <= 30'b000000010000000000011011010000
                ;mem[12647] <= 30'b000000010000000000011100100000
                ;mem[12648] <= 30'b000000010000000000011100110000
                ;mem[12649] <= 30'b000000010000000000100001100000
                ;mem[12650] <= 30'b000000010000000000100001110000
                ;mem[12651] <= 30'b000000010000000000100010000000
                ;mem[12652] <= 30'b000000010000000000100010010000
                ;mem[12653] <= 30'b000000010000000000100011100000
                ;mem[12654] <= 30'b000000010000000000100011110000
                ;mem[12655] <= 30'b000000010000000000101000100000
                ;mem[12656] <= 30'b000000010000000000101000110000
                ;mem[12657] <= 30'b000000010000000000101001000000
                ;mem[12658] <= 30'b000000010000000000101010100000
                ;mem[12659] <= 30'b000000010000000000101010110000
                ;mem[12660] <= 30'b000000010000000000101111110000
                ;mem[12661] <= 30'b000000010000000000110000000000
                ;mem[12662] <= 30'b000000010000000000110000010000
                ;mem[12663] <= 30'b000000010000000000110000100000
                ;mem[12664] <= 30'b000000010000000000110000110000
                ;mem[12665] <= 30'b000000010000000000110001000000
                ;mem[12666] <= 30'b000000010000000000110001010000
                ;mem[12667] <= 30'b000000010000000000110001100000
                ;mem[12668] <= 30'b000000010000000000110111000000
                ;mem[12669] <= 30'b000000010000000000110111010000
                ;mem[12670] <= 30'b000000010000000000110111100000
                ;mem[12671] <= 30'b000000010000000000110111110000
                ;mem[12672] <= 30'b000000010000000000111000000000
                ;mem[12673] <= 30'b000000010000000000111000010000
                ;mem[12674] <= 30'b000000010000000000111000100000
                ;mem[12675] <= 30'b000000010000000000111110010000
                ;mem[12676] <= 30'b000000010000000000111110100000
                ;mem[12677] <= 30'b000000010000000000111110110000
                ;mem[12678] <= 30'b000000010000000000111111000000
                ;mem[12679] <= 30'b000000010000000000111111010000
                ;mem[12680] <= 30'b000000000000000001000011110000
                ;mem[12681] <= 30'b000000000000000001000100000000
                ;mem[12682] <= 30'b000000000000000001000100010000
                ;mem[12683] <= 30'b000000000000000001000100100000
                ;mem[12684] <= 30'b000000000000000001000100110000
                ;mem[12685] <= 30'b000000000000000001000101000000
                ;mem[12686] <= 30'b000000000000000001000101010000
                ;mem[12687] <= 30'b000000000000000001000101100000
                ;mem[12688] <= 30'b000000000000000001001011000000
                ;mem[12689] <= 30'b000000000000000001001011010000
                ;mem[12690] <= 30'b000000000000000001001011100000
                ;mem[12691] <= 30'b000000000000000001001011110000
                ;mem[12692] <= 30'b000000000000000001001100000000
                ;mem[12693] <= 30'b000000000000000001001100010000
                ;mem[12694] <= 30'b000000000000000001001100100000
                ;mem[12695] <= 30'b000000000000000001010010010000
                ;mem[12696] <= 30'b000000000000000001010010100000
                ;mem[12697] <= 30'b000000000000000001010010110000
                ;mem[12698] <= 30'b000000000000000001010011000000
                ;mem[12699] <= 30'b000000000000000001010011010000
                ;mem[12700] <= 30'b000000000000000000101110000000
                ;mem[12701] <= 30'b000000000000000000101110010000
                ;mem[12702] <= 30'b000000000000000000101110100000
                ;mem[12703] <= 30'b000000000000000000110100100000
                ;mem[12704] <= 30'b000000000000000000110100110000
                ;mem[12705] <= 30'b000000000000000000110101100000
                ;mem[12706] <= 30'b000000000000000000110110010000
                ;mem[12707] <= 30'b000000000000000000110110100000
                ;mem[12708] <= 30'b000000000000000000111011010000
                ;mem[12709] <= 30'b000000000000000000111011100000
                ;mem[12710] <= 30'b000000000000000000111101000000
                ;mem[12711] <= 30'b000000000000000000111101010000
                ;mem[12712] <= 30'b000000001000000000000010000000
                ;mem[12713] <= 30'b000000001000000000000010010000
                ;mem[12714] <= 30'b000000001000000000000010100000
                ;mem[12715] <= 30'b000000001000000000001000100000
                ;mem[12716] <= 30'b000000001000000000001000110000
                ;mem[12717] <= 30'b000000001000000000001001100000
                ;mem[12718] <= 30'b000000001000000000001010010000
                ;mem[12719] <= 30'b000000001000000000001010100000
                ;mem[12720] <= 30'b000000001000000000001111010000
                ;mem[12721] <= 30'b000000001000000000001111100000
                ;mem[12722] <= 30'b000000001000000000010001000000
                ;mem[12723] <= 30'b000000001000000000010001010000
                ;mem[12724] <= 30'b000000001000000000010110010000
                ;mem[12725] <= 30'b000000001000000000011000000000
                ;mem[12726] <= 30'b000000001000000000011101010000
                ;mem[12727] <= 30'b000000001000000000011110110000
                ;mem[12728] <= 30'b000000001000000000011111000000
                ;mem[12729] <= 30'b000000001000000000100011110000
                ;mem[12730] <= 30'b000000001000000000100100000000
                ;mem[12731] <= 30'b000000001000000000100101100000
                ;mem[12732] <= 30'b000000001000000000100101110000
                ;mem[12733] <= 30'b000000001000000000101010110000
                ;mem[12734] <= 30'b000000001000000000101100010000
                ;mem[12735] <= 30'b000000001000000000101100100000
                ;mem[12736] <= 30'b000000001000000000101100110000
                ;mem[12737] <= 30'b000000001000000000110001100000
                ;mem[12738] <= 30'b000000001000000000110011000000
                ;mem[12739] <= 30'b000000001000000000110011010000
                ;mem[12740] <= 30'b000000001000000000111000100000
                ;mem[12741] <= 30'b000000001000000000111001100000
                ;mem[12742] <= 30'b000000001000000000111001110000
                ;mem[12743] <= 30'b000000001000000000111010000000
                ;mem[12744] <= 30'b000000001000000000111111100000
                ;mem[12745] <= 30'b000000001000000000111111110000
                ;mem[12746] <= 30'b000000010000000000000000010000
                ;mem[12747] <= 30'b000000010000000000000000100000
                ;mem[12748] <= 30'b000000010000000000000000110000
                ;mem[12749] <= 30'b000000010000000000000101100000
                ;mem[12750] <= 30'b000000010000000000000111000000
                ;mem[12751] <= 30'b000000010000000000000111010000
                ;mem[12752] <= 30'b000000010000000000001100100000
                ;mem[12753] <= 30'b000000010000000000001101100000
                ;mem[12754] <= 30'b000000010000000000001101110000
                ;mem[12755] <= 30'b000000010000000000001110000000
                ;mem[12756] <= 30'b000000010000000000010011100000
                ;mem[12757] <= 30'b000000010000000000010011110000
                ;mem[12758] <= 30'b000000010000000000010100000000
                ;mem[12759] <= 30'b000000010000000000010100010000
                ;mem[12760] <= 30'b000000010000000000010100100000
                ;mem[12761] <= 30'b000000010000000000010100110000
                ;mem[12762] <= 30'b000000010000000000010101000000
                ;mem[12763] <= 30'b000000010000000000011010110000
                ;mem[12764] <= 30'b000000010000000000011011100000
                ;mem[12765] <= 30'b000000010000000000011011110000
                ;mem[12766] <= 30'b000000010000000000011100000000
                ;mem[12767] <= 30'b000000010000000000100010100000
                ;mem[12768] <= 30'b000000010000000000100010110000
                ;mem[12769] <= 30'b000000010000000000101001010000
                ;mem[12770] <= 30'b000000010000000000101001100000
                ;mem[12771] <= 30'b000000010000000000110000000000
                ;mem[12772] <= 30'b000000010000000000110000010000
                ;mem[12773] <= 30'b000000010000000000110111000000
                ;mem[12774] <= 30'b000000010000000000111101110000
                ;mem[12775] <= 30'b000000000000000001000100000000
                ;mem[12776] <= 30'b000000000000000001000100010000
                ;mem[12777] <= 30'b000000000000000001001011000000
                ;mem[12778] <= 30'b000000000000000001010001110000
                ;mem[12779] <= 30'b000000000000000001011000100000
                ;mem[12780] <= 30'b000000000000000001011000110000
                ;mem[12781] <= 30'b000000000000000001011111010000
                ;mem[12782] <= 30'b000000000000000001011111100000
                ;mem[12783] <= 30'b000000000000000001100110010000
                ;mem[12784] <= 30'b000000000000000000100110010000
                ;mem[12785] <= 30'b000000000000000000100110100000
                ;mem[12786] <= 30'b000000000000000000101100000000
                ;mem[12787] <= 30'b000000000000000000101100010000
                ;mem[12788] <= 30'b000000000000000000101100100000
                ;mem[12789] <= 30'b000000000000000000101100110000
                ;mem[12790] <= 30'b000000000000000000101101000000
                ;mem[12791] <= 30'b000000000000000000101101010000
                ;mem[12792] <= 30'b000000000000000000101101100000
                ;mem[12793] <= 30'b000000000000000000101101110000
                ;mem[12794] <= 30'b000000000000000000101110000000
                ;mem[12795] <= 30'b000000000000000000110011000000
                ;mem[12796] <= 30'b000000000000000000110011010000
                ;mem[12797] <= 30'b000000000000000000110011100000
                ;mem[12798] <= 30'b000000000000000000110011110000
                ;mem[12799] <= 30'b000000000000000000110100000000
                ;mem[12800] <= 30'b000000000000000000110100010000
                ;mem[12801] <= 30'b000000000000000000110100100000
                ;mem[12802] <= 30'b000000000000000000110100110000
                ;mem[12803] <= 30'b000000000000000000110101000000
                ;mem[12804] <= 30'b000000000000000000110101010000
                ;mem[12805] <= 30'b000000000000000000110101100000
                ;mem[12806] <= 30'b000000000000000000111010100000
                ;mem[12807] <= 30'b000000000000000000111010110000
                ;mem[12808] <= 30'b000000000000000000111011000000
                ;mem[12809] <= 30'b000000000000000000111011010000
                ;mem[12810] <= 30'b000000000000000000111011100000
                ;mem[12811] <= 30'b000000000000000000111011110000
                ;mem[12812] <= 30'b000000000000000000111100000000
                ;mem[12813] <= 30'b000000000000000000111100010000
                ;mem[12814] <= 30'b000000000000000000111100100000
                ;mem[12815] <= 30'b000000001000000000000000000000
                ;mem[12816] <= 30'b000000001000000000000000010000
                ;mem[12817] <= 30'b000000001000000000000000100000
                ;mem[12818] <= 30'b000000001000000000000000110000
                ;mem[12819] <= 30'b000000001000000000000001000000
                ;mem[12820] <= 30'b000000001000000000000001010000
                ;mem[12821] <= 30'b000000001000000000000001100000
                ;mem[12822] <= 30'b000000001000000000000001110000
                ;mem[12823] <= 30'b000000001000000000000010000000
                ;mem[12824] <= 30'b000000001000000000000111000000
                ;mem[12825] <= 30'b000000001000000000000111010000
                ;mem[12826] <= 30'b000000001000000000000111100000
                ;mem[12827] <= 30'b000000001000000000000111110000
                ;mem[12828] <= 30'b000000001000000000001000000000
                ;mem[12829] <= 30'b000000001000000000001000010000
                ;mem[12830] <= 30'b000000001000000000001000100000
                ;mem[12831] <= 30'b000000001000000000001000110000
                ;mem[12832] <= 30'b000000001000000000001001000000
                ;mem[12833] <= 30'b000000001000000000001001010000
                ;mem[12834] <= 30'b000000001000000000001001100000
                ;mem[12835] <= 30'b000000001000000000001110100000
                ;mem[12836] <= 30'b000000001000000000001110110000
                ;mem[12837] <= 30'b000000001000000000001111000000
                ;mem[12838] <= 30'b000000001000000000001111010000
                ;mem[12839] <= 30'b000000001000000000001111100000
                ;mem[12840] <= 30'b000000001000000000001111110000
                ;mem[12841] <= 30'b000000001000000000010000000000
                ;mem[12842] <= 30'b000000001000000000010000010000
                ;mem[12843] <= 30'b000000001000000000010000100000
                ;mem[12844] <= 30'b000000001000000000010101110000
                ;mem[12845] <= 30'b000000001000000000010110000000
                ;mem[12846] <= 30'b000000001000000000010110010000
                ;mem[12847] <= 30'b000000001000000000010110100000
                ;mem[12848] <= 30'b000000001000000000010110110000
                ;mem[12849] <= 30'b000000001000000000010111000000
                ;mem[12850] <= 30'b000000001000000000010111010000
                ;mem[12851] <= 30'b000000001000000000010111100000
                ;mem[12852] <= 30'b000000001000000000011100110000
                ;mem[12853] <= 30'b000000001000000000011101000000
                ;mem[12854] <= 30'b000000001000000000011101010000
                ;mem[12855] <= 30'b000000001000000000011101100000
                ;mem[12856] <= 30'b000000001000000000011101110000
                ;mem[12857] <= 30'b000000001000000000011110000000
                ;mem[12858] <= 30'b000000001000000000011110010000
                ;mem[12859] <= 30'b000000001000000000011110100000
                ;mem[12860] <= 30'b000000001000000000100011110000
                ;mem[12861] <= 30'b000000001000000000100100000000
                ;mem[12862] <= 30'b000000001000000000100100010000
                ;mem[12863] <= 30'b000000001000000000100100100000
                ;mem[12864] <= 30'b000000001000000000100100110000
                ;mem[12865] <= 30'b000000001000000000100101000000
                ;mem[12866] <= 30'b000000001000000000100101010000
                ;mem[12867] <= 30'b000000001000000000101010100000
                ;mem[12868] <= 30'b000000001000000000101010110000
                ;mem[12869] <= 30'b000000001000000000101011000000
                ;mem[12870] <= 30'b000000001000000000101011010000
                ;mem[12871] <= 30'b000000001000000000101011100000
                ;mem[12872] <= 30'b000000001000000000101011110000
                ;mem[12873] <= 30'b000000001000000000101100000000
                ;mem[12874] <= 30'b000000001000000000101100010000
                ;mem[12875] <= 30'b000000001000000000101100100000
                ;mem[12876] <= 30'b000000001000000000110001110000
                ;mem[12877] <= 30'b000000001000000000110010000000
                ;mem[12878] <= 30'b000000001000000000110010010000
                ;mem[12879] <= 30'b000000001000000000110010100000
                ;mem[12880] <= 30'b000000001000000000110010110000
                ;mem[12881] <= 30'b000000001000000000110011000000
                ;mem[12882] <= 30'b000000001000000000110011010000
                ;mem[12883] <= 30'b000000001000000000110011100000
                ;mem[12884] <= 30'b000000001000000000111001000000
                ;mem[12885] <= 30'b000000001000000000111001010000
                ;mem[12886] <= 30'b000000001000000000111001100000
                ;mem[12887] <= 30'b000000001000000000111001110000
                ;mem[12888] <= 30'b000000001000000000111010000000
                ;mem[12889] <= 30'b000000001000000000111010010000
                ;mem[12890] <= 30'b000000001000000000111010100000
                ;mem[12891] <= 30'b000000010000000000000000000000
                ;mem[12892] <= 30'b000000010000000000000000010000
                ;mem[12893] <= 30'b000000010000000000000000100000
                ;mem[12894] <= 30'b000000010000000000000101110000
                ;mem[12895] <= 30'b000000010000000000000110000000
                ;mem[12896] <= 30'b000000010000000000000110010000
                ;mem[12897] <= 30'b000000010000000000000110100000
                ;mem[12898] <= 30'b000000010000000000000110110000
                ;mem[12899] <= 30'b000000010000000000000111000000
                ;mem[12900] <= 30'b000000010000000000000111010000
                ;mem[12901] <= 30'b000000010000000000000111100000
                ;mem[12902] <= 30'b000000010000000000001101000000
                ;mem[12903] <= 30'b000000010000000000001101010000
                ;mem[12904] <= 30'b000000010000000000001101100000
                ;mem[12905] <= 30'b000000010000000000001101110000
                ;mem[12906] <= 30'b000000010000000000001110000000
                ;mem[12907] <= 30'b000000010000000000001110010000
                ;mem[12908] <= 30'b000000010000000000001110100000
                ;mem[12909] <= 30'b000000010000000000010100110000
                ;mem[12910] <= 30'b000000010000000000010101000000
                ;mem[12911] <= 30'b000000010000000000010101010000
                ;mem[12912] <= 30'b000000010000000000010101100000
                ;mem[12913] <= 30'b000000010000000000010101110000
                ;mem[12914] <= 30'b000000010000000000011100000000
                ;mem[12915] <= 30'b000000010000000000011100010000
                ;mem[12916] <= 30'b000000010000000000011100100000
                ;mem[12917] <= 30'b000000010000000000011100110000
                ;mem[12918] <= 30'b000000010000000000100011000000
                ;mem[12919] <= 30'b000000010000000000100011010000
                ;mem[12920] <= 30'b000000010000000000100011100000
                ;mem[12921] <= 30'b000000010000000000100011110000
                ;mem[12922] <= 30'b000000010000000000101001110000
                ;mem[12923] <= 30'b000000010000000000101010000000
                ;mem[12924] <= 30'b000000010000000000101010010000
                ;mem[12925] <= 30'b000000010000000000101010100000
                ;mem[12926] <= 30'b000000010000000000110000100000
                ;mem[12927] <= 30'b000000010000000000110000110000
                ;mem[12928] <= 30'b000000010000000000110001000000
                ;mem[12929] <= 30'b000000010000000000110001010000
                ;mem[12930] <= 30'b000000010000000000110001100000
                ;mem[12931] <= 30'b000000010000000000110110000000
                ;mem[12932] <= 30'b000000010000000000110110010000
                ;mem[12933] <= 30'b000000010000000000110110100000
                ;mem[12934] <= 30'b000000010000000000110111000000
                ;mem[12935] <= 30'b000000010000000000110111010000
                ;mem[12936] <= 30'b000000010000000000110111100000
                ;mem[12937] <= 30'b000000010000000000110111110000
                ;mem[12938] <= 30'b000000010000000000111000000000
                ;mem[12939] <= 30'b000000010000000000111000010000
                ;mem[12940] <= 30'b000000010000000000111000100000
                ;mem[12941] <= 30'b000000010000000000111101000000
                ;mem[12942] <= 30'b000000010000000000111101010000
                ;mem[12943] <= 30'b000000010000000000111101100000
                ;mem[12944] <= 30'b000000010000000000111101110000
                ;mem[12945] <= 30'b000000010000000000111110000000
                ;mem[12946] <= 30'b000000010000000000111110010000
                ;mem[12947] <= 30'b000000010000000000111110100000
                ;mem[12948] <= 30'b000000010000000000111110110000
                ;mem[12949] <= 30'b000000010000000000111111000000
                ;mem[12950] <= 30'b000000010000000000111111010000
                ;mem[12951] <= 30'b000000000000000001000100100000
                ;mem[12952] <= 30'b000000000000000001000100110000
                ;mem[12953] <= 30'b000000000000000001000101000000
                ;mem[12954] <= 30'b000000000000000001000101010000
                ;mem[12955] <= 30'b000000000000000001000101100000
                ;mem[12956] <= 30'b000000000000000001001010000000
                ;mem[12957] <= 30'b000000000000000001001010010000
                ;mem[12958] <= 30'b000000000000000001001010100000
                ;mem[12959] <= 30'b000000000000000001001011000000
                ;mem[12960] <= 30'b000000000000000001001011010000
                ;mem[12961] <= 30'b000000000000000001001011100000
                ;mem[12962] <= 30'b000000000000000001001011110000
                ;mem[12963] <= 30'b000000000000000001001100000000
                ;mem[12964] <= 30'b000000000000000001001100010000
                ;mem[12965] <= 30'b000000000000000001001100100000
                ;mem[12966] <= 30'b000000000000000001010001000000
                ;mem[12967] <= 30'b000000000000000001010001010000
                ;mem[12968] <= 30'b000000000000000001010001100000
                ;mem[12969] <= 30'b000000000000000001010001110000
                ;mem[12970] <= 30'b000000000000000001010010000000
                ;mem[12971] <= 30'b000000000000000001010010010000
                ;mem[12972] <= 30'b000000000000000001010010100000
                ;mem[12973] <= 30'b000000000000000001010010110000
                ;mem[12974] <= 30'b000000000000000001010011000000
                ;mem[12975] <= 30'b000000000000000001010011010000
                ;mem[12976] <= 30'b000000000000000001011000000000
                ;mem[12977] <= 30'b000000000000000001011000010000
                ;mem[12978] <= 30'b000000000000000001011000100000
                ;mem[12979] <= 30'b000000000000000001011000110000
                ;mem[12980] <= 30'b000000000000000001011001000000
                ;mem[12981] <= 30'b000000000000000001011001010000
                ;mem[12982] <= 30'b000000000000000001011001100000
                ;mem[12983] <= 30'b000000000000000001011001110000
                ;mem[12984] <= 30'b000000000000000001011010000000
                ;mem[12985] <= 30'b000000000000000001011010010000
                ;mem[12986] <= 30'b000000000000000001011111000000
                ;mem[12987] <= 30'b000000000000000001011111010000
                ;mem[12988] <= 30'b000000000000000001011111100000
                ;mem[12989] <= 30'b000000000000000001011111110000
                ;mem[12990] <= 30'b000000000000000001100000000000
                ;mem[12991] <= 30'b000000000000000001100000010000
                ;mem[12992] <= 30'b000000000000000001100000100000
                ;mem[12993] <= 30'b000000000000000001100000110000
                ;mem[12994] <= 30'b000000000000000001100110100000
                ;mem[12995] <= 30'b000000000000000001100110110000
                ;mem[12996] <= 30'b000000000000000001100111000000
                ;mem[12997] <= 30'b000000000000000001100111010000
                ;mem[12998] <= 30'b000000000000000000011111000000
                ;mem[12999] <= 30'b000000000000000000011111010000
                ;mem[13000] <= 30'b000000000000000000011111100000
                ;mem[13001] <= 30'b000000000000000000100101110000
                ;mem[13002] <= 30'b000000000000000000100110000000
                ;mem[13003] <= 30'b000000000000000000100110010000
                ;mem[13004] <= 30'b000000000000000000100110100000
                ;mem[13005] <= 30'b000000000000000000101100110000
                ;mem[13006] <= 30'b000000000000000000101101000000
                ;mem[13007] <= 30'b000000000000000000101101010000
                ;mem[13008] <= 30'b000000000000000000101101100000
                ;mem[13009] <= 30'b000000000000000000110011110000
                ;mem[13010] <= 30'b000000000000000000110100000000
                ;mem[13011] <= 30'b000000000000000000110100010000
                ;mem[13012] <= 30'b000000000000000000110100100000
                ;mem[13013] <= 30'b000000000000000000111010110000
                ;mem[13014] <= 30'b000000000000000000111011000000
                ;mem[13015] <= 30'b000000000000000000111011010000
                ;mem[13016] <= 30'b000000000000000000111011100000
                ;mem[13017] <= 30'b000000001000000000000000110000
                ;mem[13018] <= 30'b000000001000000000000001000000
                ;mem[13019] <= 30'b000000001000000000000001010000
                ;mem[13020] <= 30'b000000001000000000000001100000
                ;mem[13021] <= 30'b000000001000000000000111110000
                ;mem[13022] <= 30'b000000001000000000001000000000
                ;mem[13023] <= 30'b000000001000000000001000010000
                ;mem[13024] <= 30'b000000001000000000001000100000
                ;mem[13025] <= 30'b000000001000000000001110110000
                ;mem[13026] <= 30'b000000001000000000001111000000
                ;mem[13027] <= 30'b000000001000000000001111010000
                ;mem[13028] <= 30'b000000001000000000001111100000
                ;mem[13029] <= 30'b000000001000000000010101110000
                ;mem[13030] <= 30'b000000001000000000010110000000
                ;mem[13031] <= 30'b000000001000000000010110010000
                ;mem[13032] <= 30'b000000001000000000010110100000
                ;mem[13033] <= 30'b000000001000000000010110110000
                ;mem[13034] <= 30'b000000001000000000011100110000
                ;mem[13035] <= 30'b000000001000000000011101000000
                ;mem[13036] <= 30'b000000001000000000011101010000
                ;mem[13037] <= 30'b000000001000000000011101100000
                ;mem[13038] <= 30'b000000001000000000011101110000
                ;mem[13039] <= 30'b000000001000000000100011110000
                ;mem[13040] <= 30'b000000001000000000100100000000
                ;mem[13041] <= 30'b000000001000000000100100010000
                ;mem[13042] <= 30'b000000001000000000100100100000
                ;mem[13043] <= 30'b000000001000000000100100110000
                ;mem[13044] <= 30'b000000001000000000100101000000
                ;mem[13045] <= 30'b000000001000000000101011000000
                ;mem[13046] <= 30'b000000001000000000101011010000
                ;mem[13047] <= 30'b000000001000000000101011100000
                ;mem[13048] <= 30'b000000001000000000101011110000
                ;mem[13049] <= 30'b000000001000000000101100000000
                ;mem[13050] <= 30'b000000001000000000110010000000
                ;mem[13051] <= 30'b000000001000000000110010010000
                ;mem[13052] <= 30'b000000001000000000110010100000
                ;mem[13053] <= 30'b000000001000000000110010110000
                ;mem[13054] <= 30'b000000001000000000110011000000
                ;mem[13055] <= 30'b000000001000000000111001000000
                ;mem[13056] <= 30'b000000001000000000111001010000
                ;mem[13057] <= 30'b000000001000000000111001100000
                ;mem[13058] <= 30'b000000001000000000111001110000
                ;mem[13059] <= 30'b000000001000000000111010000000
                ;mem[13060] <= 30'b000000010000000000000000000000
                ;mem[13061] <= 30'b000000010000000000000110000000
                ;mem[13062] <= 30'b000000010000000000000110010000
                ;mem[13063] <= 30'b000000010000000000000110100000
                ;mem[13064] <= 30'b000000010000000000000110110000
                ;mem[13065] <= 30'b000000010000000000000111000000
                ;mem[13066] <= 30'b000000010000000000001101000000
                ;mem[13067] <= 30'b000000010000000000001101010000
                ;mem[13068] <= 30'b000000010000000000001101100000
                ;mem[13069] <= 30'b000000010000000000001101110000
                ;mem[13070] <= 30'b000000010000000000001110000000
                ;mem[13071] <= 30'b000000010000000000010100000000
                ;mem[13072] <= 30'b000000010000000000010100010000
                ;mem[13073] <= 30'b000000010000000000010100100000
                ;mem[13074] <= 30'b000000010000000000010100110000
                ;mem[13075] <= 30'b000000010000000000010101000000
                ;mem[13076] <= 30'b000000010000000000011011000000
                ;mem[13077] <= 30'b000000010000000000011011010000
                ;mem[13078] <= 30'b000000010000000000011011100000
                ;mem[13079] <= 30'b000000010000000000011011110000
                ;mem[13080] <= 30'b000000010000000000011100000000
                ;mem[13081] <= 30'b000000010000000000100010000000
                ;mem[13082] <= 30'b000000010000000000100010010000
                ;mem[13083] <= 30'b000000010000000000100010100000
                ;mem[13084] <= 30'b000000010000000000100010110000
                ;mem[13085] <= 30'b000000010000000000100011000000
                ;mem[13086] <= 30'b000000010000000000101001000000
                ;mem[13087] <= 30'b000000010000000000101001010000
                ;mem[13088] <= 30'b000000010000000000101001100000
                ;mem[13089] <= 30'b000000010000000000101001110000
                ;mem[13090] <= 30'b000000010000000000101010000000
                ;mem[13091] <= 30'b000000010000000000110000000000
                ;mem[13092] <= 30'b000000010000000000110000010000
                ;mem[13093] <= 30'b000000010000000000110000100000
                ;mem[13094] <= 30'b000000010000000000110000110000
                ;mem[13095] <= 30'b000000010000000000110001000000
                ;mem[13096] <= 30'b000000010000000000110111010000
                ;mem[13097] <= 30'b000000010000000000110111100000
                ;mem[13098] <= 30'b000000010000000000110111110000
                ;mem[13099] <= 30'b000000010000000000111000000000
                ;mem[13100] <= 30'b000000010000000000111110010000
                ;mem[13101] <= 30'b000000010000000000111110100000
                ;mem[13102] <= 30'b000000010000000000111110110000
                ;mem[13103] <= 30'b000000010000000000111111000000
                ;mem[13104] <= 30'b000000010000000000111111010000
                ;mem[13105] <= 30'b000000000000000001000100000000
                ;mem[13106] <= 30'b000000000000000001000100010000
                ;mem[13107] <= 30'b000000000000000001000100100000
                ;mem[13108] <= 30'b000000000000000001000100110000
                ;mem[13109] <= 30'b000000000000000001000101000000
                ;mem[13110] <= 30'b000000000000000001001011010000
                ;mem[13111] <= 30'b000000000000000001001011100000
                ;mem[13112] <= 30'b000000000000000001001011110000
                ;mem[13113] <= 30'b000000000000000001001100000000
                ;mem[13114] <= 30'b000000000000000001010010010000
                ;mem[13115] <= 30'b000000000000000001010010100000
                ;mem[13116] <= 30'b000000000000000001010010110000
                ;mem[13117] <= 30'b000000000000000001010011000000
                ;mem[13118] <= 30'b000000000000000001010011010000
                ;mem[13119] <= 30'b000000000000000001011001010000
                ;mem[13120] <= 30'b000000000000000001011001100000
                ;mem[13121] <= 30'b000000000000000001011001110000
                ;mem[13122] <= 30'b000000000000000001011010000000
                ;mem[13123] <= 30'b000000000000000001011010010000
                ;mem[13124] <= 30'b000000000000000001011010100000
                ;mem[13125] <= 30'b000000000000000001100000110000
                ;mem[13126] <= 30'b000000000000000001100001000000
                ;mem[13127] <= 30'b000000000000000001100001010000
                ;mem[13128] <= 30'b000000000000000000100111110000
                ;mem[13129] <= 30'b000000000000000000101000000000
                ;mem[13130] <= 30'b000000000000000000101000010000
                ;mem[13131] <= 30'b000000000000000000101110100000
                ;mem[13132] <= 30'b000000000000000000101110110000
                ;mem[13133] <= 30'b000000000000000000101111000000
                ;mem[13134] <= 30'b000000000000000000101111010000
                ;mem[13135] <= 30'b000000000000000000110100000000
                ;mem[13136] <= 30'b000000000000000000110100010000
                ;mem[13137] <= 30'b000000000000000000110100100000
                ;mem[13138] <= 30'b000000000000000000110101010000
                ;mem[13139] <= 30'b000000000000000000110101100000
                ;mem[13140] <= 30'b000000000000000000110101110000
                ;mem[13141] <= 30'b000000000000000000110110000000
                ;mem[13142] <= 30'b000000000000000000110110010000
                ;mem[13143] <= 30'b000000000000000000111010110000
                ;mem[13144] <= 30'b000000000000000000111011000000
                ;mem[13145] <= 30'b000000000000000000111011010000
                ;mem[13146] <= 30'b000000000000000000111100000000
                ;mem[13147] <= 30'b000000000000000000111100010000
                ;mem[13148] <= 30'b000000000000000000111100100000
                ;mem[13149] <= 30'b000000000000000000111100110000
                ;mem[13150] <= 30'b000000000000000000111101000000
                ;mem[13151] <= 30'b000000001000000000000010100000
                ;mem[13152] <= 30'b000000001000000000000010110000
                ;mem[13153] <= 30'b000000001000000000000011000000
                ;mem[13154] <= 30'b000000001000000000000011010000
                ;mem[13155] <= 30'b000000001000000000001000000000
                ;mem[13156] <= 30'b000000001000000000001000010000
                ;mem[13157] <= 30'b000000001000000000001000100000
                ;mem[13158] <= 30'b000000001000000000001001010000
                ;mem[13159] <= 30'b000000001000000000001001100000
                ;mem[13160] <= 30'b000000001000000000001001110000
                ;mem[13161] <= 30'b000000001000000000001010000000
                ;mem[13162] <= 30'b000000001000000000001010010000
                ;mem[13163] <= 30'b000000001000000000001110110000
                ;mem[13164] <= 30'b000000001000000000001111000000
                ;mem[13165] <= 30'b000000001000000000001111010000
                ;mem[13166] <= 30'b000000001000000000010000000000
                ;mem[13167] <= 30'b000000001000000000010000010000
                ;mem[13168] <= 30'b000000001000000000010000100000
                ;mem[13169] <= 30'b000000001000000000010000110000
                ;mem[13170] <= 30'b000000001000000000010001000000
                ;mem[13171] <= 30'b000000001000000000010101100000
                ;mem[13172] <= 30'b000000001000000000010101110000
                ;mem[13173] <= 30'b000000001000000000010110000000
                ;mem[13174] <= 30'b000000001000000000010110110000
                ;mem[13175] <= 30'b000000001000000000010111000000
                ;mem[13176] <= 30'b000000001000000000010111010000
                ;mem[13177] <= 30'b000000001000000000010111100000
                ;mem[13178] <= 30'b000000001000000000011100010000
                ;mem[13179] <= 30'b000000001000000000011100100000
                ;mem[13180] <= 30'b000000001000000000011100110000
                ;mem[13181] <= 30'b000000001000000000011101110000
                ;mem[13182] <= 30'b000000001000000000011110000000
                ;mem[13183] <= 30'b000000001000000000011110010000
                ;mem[13184] <= 30'b000000001000000000011110100000
                ;mem[13185] <= 30'b000000001000000000100011000000
                ;mem[13186] <= 30'b000000001000000000100011010000
                ;mem[13187] <= 30'b000000001000000000100011100000
                ;mem[13188] <= 30'b000000001000000000100011110000
                ;mem[13189] <= 30'b000000001000000000100100100000
                ;mem[13190] <= 30'b000000001000000000100100110000
                ;mem[13191] <= 30'b000000001000000000100101000000
                ;mem[13192] <= 30'b000000001000000000100101010000
                ;mem[13193] <= 30'b000000001000000000100101100000
                ;mem[13194] <= 30'b000000001000000000101001110000
                ;mem[13195] <= 30'b000000001000000000101010000000
                ;mem[13196] <= 30'b000000001000000000101010010000
                ;mem[13197] <= 30'b000000001000000000101010100000
                ;mem[13198] <= 30'b000000001000000000101011100000
                ;mem[13199] <= 30'b000000001000000000101011110000
                ;mem[13200] <= 30'b000000001000000000101100000000
                ;mem[13201] <= 30'b000000001000000000101100010000
                ;mem[13202] <= 30'b000000001000000000101101000000
                ;mem[13203] <= 30'b000000001000000000101101010000
                ;mem[13204] <= 30'b000000001000000000110000100000
                ;mem[13205] <= 30'b000000001000000000110000110000
                ;mem[13206] <= 30'b000000001000000000110001000000
                ;mem[13207] <= 30'b000000001000000000110001010000
                ;mem[13208] <= 30'b000000001000000000110010100000
                ;mem[13209] <= 30'b000000001000000000110010110000
                ;mem[13210] <= 30'b000000001000000000110011000000
                ;mem[13211] <= 30'b000000001000000000110011010000
                ;mem[13212] <= 30'b000000001000000000110011110000
                ;mem[13213] <= 30'b000000001000000000110100000000
                ;mem[13214] <= 30'b000000001000000000110100010000
                ;mem[13215] <= 30'b000000001000000000110111100000
                ;mem[13216] <= 30'b000000001000000000110111110000
                ;mem[13217] <= 30'b000000001000000000111000000000
                ;mem[13218] <= 30'b000000001000000000111000010000
                ;mem[13219] <= 30'b000000001000000000111001100000
                ;mem[13220] <= 30'b000000001000000000111001110000
                ;mem[13221] <= 30'b000000001000000000111010000000
                ;mem[13222] <= 30'b000000001000000000111010010000
                ;mem[13223] <= 30'b000000001000000000111010100000
                ;mem[13224] <= 30'b000000001000000000111010110000
                ;mem[13225] <= 30'b000000001000000000111011000000
                ;mem[13226] <= 30'b000000001000000000111011010000
                ;mem[13227] <= 30'b000000001000000000111110100000
                ;mem[13228] <= 30'b000000001000000000111110110000
                ;mem[13229] <= 30'b000000001000000000111111000000
                ;mem[13230] <= 30'b000000001000000000111111010000
                ;mem[13231] <= 30'b000000001000000000111111100000
                ;mem[13232] <= 30'b000000001000000000111111110000
                ;mem[13233] <= 30'b000000010000000000000000000000
                ;mem[13234] <= 30'b000000010000000000000000010000
                ;mem[13235] <= 30'b000000010000000000000001000000
                ;mem[13236] <= 30'b000000010000000000000001010000
                ;mem[13237] <= 30'b000000010000000000000100100000
                ;mem[13238] <= 30'b000000010000000000000100110000
                ;mem[13239] <= 30'b000000010000000000000101000000
                ;mem[13240] <= 30'b000000010000000000000101010000
                ;mem[13241] <= 30'b000000010000000000000110100000
                ;mem[13242] <= 30'b000000010000000000000110110000
                ;mem[13243] <= 30'b000000010000000000000111000000
                ;mem[13244] <= 30'b000000010000000000000111010000
                ;mem[13245] <= 30'b000000010000000000000111110000
                ;mem[13246] <= 30'b000000010000000000001000000000
                ;mem[13247] <= 30'b000000010000000000001000010000
                ;mem[13248] <= 30'b000000010000000000001011100000
                ;mem[13249] <= 30'b000000010000000000001011110000
                ;mem[13250] <= 30'b000000010000000000001100000000
                ;mem[13251] <= 30'b000000010000000000001100010000
                ;mem[13252] <= 30'b000000010000000000001101100000
                ;mem[13253] <= 30'b000000010000000000001101110000
                ;mem[13254] <= 30'b000000010000000000001110000000
                ;mem[13255] <= 30'b000000010000000000001110010000
                ;mem[13256] <= 30'b000000010000000000001110100000
                ;mem[13257] <= 30'b000000010000000000001110110000
                ;mem[13258] <= 30'b000000010000000000001111000000
                ;mem[13259] <= 30'b000000010000000000001111010000
                ;mem[13260] <= 30'b000000010000000000010010100000
                ;mem[13261] <= 30'b000000010000000000010010110000
                ;mem[13262] <= 30'b000000010000000000010011000000
                ;mem[13263] <= 30'b000000010000000000010011010000
                ;mem[13264] <= 30'b000000010000000000010011100000
                ;mem[13265] <= 30'b000000010000000000010011110000
                ;mem[13266] <= 30'b000000010000000000010100000000
                ;mem[13267] <= 30'b000000010000000000010100010000
                ;mem[13268] <= 30'b000000010000000000010100100000
                ;mem[13269] <= 30'b000000010000000000010100110000
                ;mem[13270] <= 30'b000000010000000000010101000000
                ;mem[13271] <= 30'b000000010000000000010101010000
                ;mem[13272] <= 30'b000000010000000000010101100000
                ;mem[13273] <= 30'b000000010000000000010101110000
                ;mem[13274] <= 30'b000000010000000000010110000000
                ;mem[13275] <= 30'b000000010000000000010110010000
                ;mem[13276] <= 30'b000000010000000000011001100000
                ;mem[13277] <= 30'b000000010000000000011001110000
                ;mem[13278] <= 30'b000000010000000000011010000000
                ;mem[13279] <= 30'b000000010000000000011010010000
                ;mem[13280] <= 30'b000000010000000000011010100000
                ;mem[13281] <= 30'b000000010000000000011010110000
                ;mem[13282] <= 30'b000000010000000000011011000000
                ;mem[13283] <= 30'b000000010000000000011011010000
                ;mem[13284] <= 30'b000000010000000000011011100000
                ;mem[13285] <= 30'b000000010000000000011011110000
                ;mem[13286] <= 30'b000000010000000000011100000000
                ;mem[13287] <= 30'b000000010000000000011100010000
                ;mem[13288] <= 30'b000000010000000000011100100000
                ;mem[13289] <= 30'b000000010000000000011100110000
                ;mem[13290] <= 30'b000000010000000000011101000000
                ;mem[13291] <= 30'b000000010000000000100000100000
                ;mem[13292] <= 30'b000000010000000000100000110000
                ;mem[13293] <= 30'b000000010000000000100001000000
                ;mem[13294] <= 30'b000000010000000000100001010000
                ;mem[13295] <= 30'b000000010000000000100001100000
                ;mem[13296] <= 30'b000000010000000000100001110000
                ;mem[13297] <= 30'b000000010000000000100010000000
                ;mem[13298] <= 30'b000000010000000000100010010000
                ;mem[13299] <= 30'b000000010000000000100010100000
                ;mem[13300] <= 30'b000000010000000000100010110000
                ;mem[13301] <= 30'b000000010000000000100011000000
                ;mem[13302] <= 30'b000000010000000000100011010000
                ;mem[13303] <= 30'b000000010000000000100011100000
                ;mem[13304] <= 30'b000000010000000000100011110000
                ;mem[13305] <= 30'b000000010000000000101000000000
                ;mem[13306] <= 30'b000000010000000000101000010000
                ;mem[13307] <= 30'b000000010000000000101000100000
                ;mem[13308] <= 30'b000000010000000000101000110000
                ;mem[13309] <= 30'b000000010000000000101001000000
                ;mem[13310] <= 30'b000000010000000000101001010000
                ;mem[13311] <= 30'b000000010000000000101001100000
                ;mem[13312] <= 30'b000000010000000000101001110000
                ;mem[13313] <= 30'b000000010000000000101010000000
                ;mem[13314] <= 30'b000000010000000000101010010000
                ;mem[13315] <= 30'b000000010000000000101111110000
                ;mem[13316] <= 30'b000000010000000000110000000000
                ;mem[13317] <= 30'b000000010000000000110000010000
                ;mem[13318] <= 30'b000000010000000000110000100000
                ;mem[13319] <= 30'b000000010000000000110000110000
                ;mem[13320] <= 30'b000000010000000000110001000000
                ;mem[13321] <= 30'b000000010000000000110111000000
                ;mem[13322] <= 30'b000000010000000000110111010000
                ;mem[13323] <= 30'b000000010000000000110111100000
                ;mem[13324] <= 30'b000000010000000000110111110000
                ;mem[13325] <= 30'b000000010000000000111000000000
                ;mem[13326] <= 30'b000000010000000000111110000000
                ;mem[13327] <= 30'b000000010000000000111110010000
                ;mem[13328] <= 30'b000000010000000000111110100000
                ;mem[13329] <= 30'b000000010000000000111110110000
                ;mem[13330] <= 30'b000000010000000000111111000000
                ;mem[13331] <= 30'b000000010000000000111111010000
                ;mem[13332] <= 30'b000000010000000000111111100000
                ;mem[13333] <= 30'b000000000000000001000011110000
                ;mem[13334] <= 30'b000000000000000001000100000000
                ;mem[13335] <= 30'b000000000000000001000100010000
                ;mem[13336] <= 30'b000000000000000001000100100000
                ;mem[13337] <= 30'b000000000000000001000100110000
                ;mem[13338] <= 30'b000000000000000001000101000000
                ;mem[13339] <= 30'b000000000000000001001011000000
                ;mem[13340] <= 30'b000000000000000001001011010000
                ;mem[13341] <= 30'b000000000000000001001011100000
                ;mem[13342] <= 30'b000000000000000001001011110000
                ;mem[13343] <= 30'b000000000000000001001100000000
                ;mem[13344] <= 30'b000000000000000001010010000000
                ;mem[13345] <= 30'b000000000000000001010010010000
                ;mem[13346] <= 30'b000000000000000001010010100000
                ;mem[13347] <= 30'b000000000000000001010010110000
                ;mem[13348] <= 30'b000000000000000001010011000000
                ;mem[13349] <= 30'b000000000000000001010011010000
                ;mem[13350] <= 30'b000000000000000001010011100000
                ;mem[13351] <= 30'b000000000000000001011001010000
                ;mem[13352] <= 30'b000000000000000001011001100000
                ;mem[13353] <= 30'b000000000000000001011001110000
                ;mem[13354] <= 30'b000000000000000001011010000000
                ;mem[13355] <= 30'b000000000000000001011010010000
                ;mem[13356] <= 30'b000000000000000001011010100000
                ;mem[13357] <= 30'b000000000000000001100000100000
                ;mem[13358] <= 30'b000000000000000001100000110000
                ;mem[13359] <= 30'b000000000000000001100001000000
                ;mem[13360] <= 30'b000000000000000001100001010000
                ;mem[13361] <= 30'b000000000000000001100111110000
                ;mem[13362] <= 30'b000000000000000000100101100000
                ;mem[13363] <= 30'b000000000000000000101100110000
                ;mem[13364] <= 30'b000000000000000000101101000000
                ;mem[13365] <= 30'b000000000000000000101101010000
                ;mem[13366] <= 30'b000000000000000000110011110000
                ;mem[13367] <= 30'b000000000000000000110100000000
                ;mem[13368] <= 30'b000000000000000000110100010000
                ;mem[13369] <= 30'b000000000000000000111010110000
                ;mem[13370] <= 30'b000000000000000000111011000000
                ;mem[13371] <= 30'b000000000000000000111011010000
                ;mem[13372] <= 30'b000000001000000000000000110000
                ;mem[13373] <= 30'b000000001000000000000001000000
                ;mem[13374] <= 30'b000000001000000000000001010000
                ;mem[13375] <= 30'b000000001000000000000111110000
                ;mem[13376] <= 30'b000000001000000000001000000000
                ;mem[13377] <= 30'b000000001000000000001000010000
                ;mem[13378] <= 30'b000000001000000000001110110000
                ;mem[13379] <= 30'b000000001000000000001111000000
                ;mem[13380] <= 30'b000000001000000000001111010000
                ;mem[13381] <= 30'b000000001000000000010101110000
                ;mem[13382] <= 30'b000000001000000000010110000000
                ;mem[13383] <= 30'b000000001000000000010110010000
                ;mem[13384] <= 30'b000000001000000000011101000000
                ;mem[13385] <= 30'b000000001000000000011101010000
                ;mem[13386] <= 30'b000000001000000000011101100000
                ;mem[13387] <= 30'b000000001000000000100100000000
                ;mem[13388] <= 30'b000000001000000000100100010000
                ;mem[13389] <= 30'b000000001000000000100100100000
                ;mem[13390] <= 30'b000000001000000000101011010000
                ;mem[13391] <= 30'b000000001000000000101011100000
                ;mem[13392] <= 30'b000000001000000000101011110000
                ;mem[13393] <= 30'b000000001000000000110010100000
                ;mem[13394] <= 30'b000000001000000000110010110000
                ;mem[13395] <= 30'b000000001000000000111001100000
                ;mem[13396] <= 30'b000000001000000000111001110000
                ;mem[13397] <= 30'b000000001000000000111010000000
                ;mem[13398] <= 30'b000000010000000000000110100000
                ;mem[13399] <= 30'b000000010000000000000110110000
                ;mem[13400] <= 30'b000000010000000000001101100000
                ;mem[13401] <= 30'b000000010000000000001101110000
                ;mem[13402] <= 30'b000000010000000000001110000000
                ;mem[13403] <= 30'b000000010000000000010100100000
                ;mem[13404] <= 30'b000000010000000000010100110000
                ;mem[13405] <= 30'b000000010000000000010101000000
                ;mem[13406] <= 30'b000000010000000000011011100000
                ;mem[13407] <= 30'b000000010000000000011011110000
                ;mem[13408] <= 30'b000000010000000000011100000000
                ;mem[13409] <= 30'b000000010000000000100010110000
                ;mem[13410] <= 30'b000000010000000000100011000000
                ;mem[13411] <= 30'b000000010000000000101001110000
                ;mem[13412] <= 30'b000000010000000000101010000000
                ;mem[13413] <= 30'b000000010000000000110001000000
                ;mem[13414] <= 30'b000000010000000000110001010000
                ;mem[13415] <= 30'b000000010000000000111000000000
                ;mem[13416] <= 30'b000000010000000000111000010000
                ;mem[13417] <= 30'b000000010000000000111111000000
                ;mem[13418] <= 30'b000000010000000000111111010000
                ;mem[13419] <= 30'b000000000000000001000101000000
                ;mem[13420] <= 30'b000000000000000001000101010000
                ;mem[13421] <= 30'b000000000000000001001100000000
                ;mem[13422] <= 30'b000000000000000001001100010000
                ;mem[13423] <= 30'b000000000000000001010011000000
                ;mem[13424] <= 30'b000000000000000001010011010000
                ;mem[13425] <= 30'b000000000000000001011010000000
                ;mem[13426] <= 30'b000000000000000001011010010000
                ;mem[13427] <= 30'b000000000000000001100001000000
                ;mem[13428] <= 30'b000000000000000001100001010000
                ;mem[13429] <= 30'b000000000000000001101000000000
                ;mem[13430] <= 30'b000000000000000000101100000000
                ;mem[13431] <= 30'b000000000000000000101110000000
                ;mem[13432] <= 30'b000000000000000000110010110000
                ;mem[13433] <= 30'b000000000000000000110011000000
                ;mem[13434] <= 30'b000000000000000000110011010000
                ;mem[13435] <= 30'b000000000000000000110011100000
                ;mem[13436] <= 30'b000000000000000000110011110000
                ;mem[13437] <= 30'b000000000000000000110100000000
                ;mem[13438] <= 30'b000000000000000000110100010000
                ;mem[13439] <= 30'b000000000000000000110100100000
                ;mem[13440] <= 30'b000000000000000000110100110000
                ;mem[13441] <= 30'b000000000000000000110101000000
                ;mem[13442] <= 30'b000000000000000000110101010000
                ;mem[13443] <= 30'b000000000000000000111001110000
                ;mem[13444] <= 30'b000000000000000000111010000000
                ;mem[13445] <= 30'b000000000000000000111010010000
                ;mem[13446] <= 30'b000000000000000000111010100000
                ;mem[13447] <= 30'b000000000000000000111010110000
                ;mem[13448] <= 30'b000000000000000000111011000000
                ;mem[13449] <= 30'b000000000000000000111011010000
                ;mem[13450] <= 30'b000000000000000000111011100000
                ;mem[13451] <= 30'b000000000000000000111011110000
                ;mem[13452] <= 30'b000000000000000000111100000000
                ;mem[13453] <= 30'b000000000000000000111100010000
                ;mem[13454] <= 30'b000000001000000000000000000000
                ;mem[13455] <= 30'b000000001000000000000010000000
                ;mem[13456] <= 30'b000000001000000000000110110000
                ;mem[13457] <= 30'b000000001000000000000111000000
                ;mem[13458] <= 30'b000000001000000000000111010000
                ;mem[13459] <= 30'b000000001000000000000111100000
                ;mem[13460] <= 30'b000000001000000000000111110000
                ;mem[13461] <= 30'b000000001000000000001000000000
                ;mem[13462] <= 30'b000000001000000000001000010000
                ;mem[13463] <= 30'b000000001000000000001000100000
                ;mem[13464] <= 30'b000000001000000000001000110000
                ;mem[13465] <= 30'b000000001000000000001001000000
                ;mem[13466] <= 30'b000000001000000000001001010000
                ;mem[13467] <= 30'b000000001000000000001101110000
                ;mem[13468] <= 30'b000000001000000000001110000000
                ;mem[13469] <= 30'b000000001000000000001110010000
                ;mem[13470] <= 30'b000000001000000000001110100000
                ;mem[13471] <= 30'b000000001000000000001110110000
                ;mem[13472] <= 30'b000000001000000000001111000000
                ;mem[13473] <= 30'b000000001000000000001111010000
                ;mem[13474] <= 30'b000000001000000000001111100000
                ;mem[13475] <= 30'b000000001000000000001111110000
                ;mem[13476] <= 30'b000000001000000000010000000000
                ;mem[13477] <= 30'b000000001000000000010000010000
                ;mem[13478] <= 30'b000000001000000000010101000000
                ;mem[13479] <= 30'b000000001000000000010101010000
                ;mem[13480] <= 30'b000000001000000000010101110000
                ;mem[13481] <= 30'b000000001000000000010110000000
                ;mem[13482] <= 30'b000000001000000000010110010000
                ;mem[13483] <= 30'b000000001000000000010110100000
                ;mem[13484] <= 30'b000000001000000000010110110000
                ;mem[13485] <= 30'b000000001000000000010111000000
                ;mem[13486] <= 30'b000000001000000000010111010000
                ;mem[13487] <= 30'b000000001000000000011101010000
                ;mem[13488] <= 30'b000000001000000000011101100000
                ;mem[13489] <= 30'b000000001000000000011101110000
                ;mem[13490] <= 30'b000000001000000000011110000000
                ;mem[13491] <= 30'b000000001000000000100100010000
                ;mem[13492] <= 30'b000000001000000000100100100000
                ;mem[13493] <= 30'b000000001000000000100100110000
                ;mem[13494] <= 30'b000000001000000000100101000000
                ;mem[13495] <= 30'b000000001000000000101011010000
                ;mem[13496] <= 30'b000000001000000000101011100000
                ;mem[13497] <= 30'b000000001000000000101011110000
                ;mem[13498] <= 30'b000000001000000000101100000000
                ;mem[13499] <= 30'b000000001000000000110001110000
                ;mem[13500] <= 30'b000000001000000000110010000000
                ;mem[13501] <= 30'b000000001000000000110010010000
                ;mem[13502] <= 30'b000000001000000000110010100000
                ;mem[13503] <= 30'b000000001000000000110010110000
                ;mem[13504] <= 30'b000000001000000000111000010000
                ;mem[13505] <= 30'b000000001000000000111000100000
                ;mem[13506] <= 30'b000000001000000000111000110000
                ;mem[13507] <= 30'b000000001000000000111001000000
                ;mem[13508] <= 30'b000000001000000000111001010000
                ;mem[13509] <= 30'b000000001000000000111001100000
                ;mem[13510] <= 30'b000000001000000000111001110000
                ;mem[13511] <= 30'b000000001000000000111010000000
                ;mem[13512] <= 30'b000000001000000000111010010000
                ;mem[13513] <= 30'b000000001000000000111010100000
                ;mem[13514] <= 30'b000000001000000000111010110000
                ;mem[13515] <= 30'b000000001000000000111011000000
                ;mem[13516] <= 30'b000000001000000000111011010000
                ;mem[13517] <= 30'b000000001000000000111011100000
                ;mem[13518] <= 30'b000000001000000000111011110000
                ;mem[13519] <= 30'b000000001000000000111100000000
                ;mem[13520] <= 30'b000000001000000000111100010000
                ;mem[13521] <= 30'b000000001000000000111100100000
                ;mem[13522] <= 30'b000000001000000000111111110000
                ;mem[13523] <= 30'b000000010000000000000000000000
                ;mem[13524] <= 30'b000000010000000000000101110000
                ;mem[13525] <= 30'b000000010000000000000110000000
                ;mem[13526] <= 30'b000000010000000000000110010000
                ;mem[13527] <= 30'b000000010000000000000110100000
                ;mem[13528] <= 30'b000000010000000000000110110000
                ;mem[13529] <= 30'b000000010000000000001100010000
                ;mem[13530] <= 30'b000000010000000000001100100000
                ;mem[13531] <= 30'b000000010000000000001100110000
                ;mem[13532] <= 30'b000000010000000000001101000000
                ;mem[13533] <= 30'b000000010000000000001101010000
                ;mem[13534] <= 30'b000000010000000000001101100000
                ;mem[13535] <= 30'b000000010000000000001101110000
                ;mem[13536] <= 30'b000000010000000000001110000000
                ;mem[13537] <= 30'b000000010000000000001110010000
                ;mem[13538] <= 30'b000000010000000000001110100000
                ;mem[13539] <= 30'b000000010000000000001110110000
                ;mem[13540] <= 30'b000000010000000000001111000000
                ;mem[13541] <= 30'b000000010000000000001111010000
                ;mem[13542] <= 30'b000000010000000000001111100000
                ;mem[13543] <= 30'b000000010000000000001111110000
                ;mem[13544] <= 30'b000000010000000000010000000000
                ;mem[13545] <= 30'b000000010000000000010000010000
                ;mem[13546] <= 30'b000000010000000000010000100000
                ;mem[13547] <= 30'b000000010000000000010011110000
                ;mem[13548] <= 30'b000000010000000000010100000000
                ;mem[13549] <= 30'b000000010000000000010100010000
                ;mem[13550] <= 30'b000000010000000000010100100000
                ;mem[13551] <= 30'b000000010000000000010100110000
                ;mem[13552] <= 30'b000000010000000000010101000000
                ;mem[13553] <= 30'b000000010000000000010101010000
                ;mem[13554] <= 30'b000000010000000000010101100000
                ;mem[13555] <= 30'b000000010000000000010101110000
                ;mem[13556] <= 30'b000000010000000000010110000000
                ;mem[13557] <= 30'b000000010000000000010110010000
                ;mem[13558] <= 30'b000000010000000000010110100000
                ;mem[13559] <= 30'b000000010000000000010110110000
                ;mem[13560] <= 30'b000000010000000000010111000000
                ;mem[13561] <= 30'b000000010000000000011011000000
                ;mem[13562] <= 30'b000000010000000000011011010000
                ;mem[13563] <= 30'b000000010000000000011011100000
                ;mem[13564] <= 30'b000000010000000000011011110000
                ;mem[13565] <= 30'b000000010000000000011100000000
                ;mem[13566] <= 30'b000000010000000000011100010000
                ;mem[13567] <= 30'b000000010000000000011100100000
                ;mem[13568] <= 30'b000000010000000000100010000000
                ;mem[13569] <= 30'b000000010000000000100010010000
                ;mem[13570] <= 30'b000000010000000000100010100000
                ;mem[13571] <= 30'b000000010000000000100010110000
                ;mem[13572] <= 30'b000000010000000000101001000000
                ;mem[13573] <= 30'b000000010000000000101001010000
                ;mem[13574] <= 30'b000000010000000000101001100000
                ;mem[13575] <= 30'b000000010000000000110000000000
                ;mem[13576] <= 30'b000000010000000000110000010000
                ;mem[13577] <= 30'b000000010000000000110000100000
                ;mem[13578] <= 30'b000000010000000000110111000000
                ;mem[13579] <= 30'b000000010000000000110111010000
                ;mem[13580] <= 30'b000000010000000000110111100000
                ;mem[13581] <= 30'b000000010000000000111110000000
                ;mem[13582] <= 30'b000000010000000000111110010000
                ;mem[13583] <= 30'b000000010000000000111110100000
                ;mem[13584] <= 30'b000000000000000001000100000000
                ;mem[13585] <= 30'b000000000000000001000100010000
                ;mem[13586] <= 30'b000000000000000001000100100000
                ;mem[13587] <= 30'b000000000000000001001011000000
                ;mem[13588] <= 30'b000000000000000001001011010000
                ;mem[13589] <= 30'b000000000000000001001011100000
                ;mem[13590] <= 30'b000000000000000001010010000000
                ;mem[13591] <= 30'b000000000000000001010010010000
                ;mem[13592] <= 30'b000000000000000001010010100000
                ;mem[13593] <= 30'b000000000000000001011001000000
                ;mem[13594] <= 30'b000000000000000001011001010000
                ;mem[13595] <= 30'b000000000000000001011001100000
                ;mem[13596] <= 30'b000000000000000001100000000000
                ;mem[13597] <= 30'b000000000000000001100000010000
                ;mem[13598] <= 30'b000000000000000001100000100000
                ;mem[13599] <= 30'b000000000000000001100111000000
                ;mem[13600] <= 30'b000000000000000001100111010000
                ;mem[13601] <= 30'b000000000000000001100111100000
                ;mem[13602] <= 30'b000000000000000001101110010000
                ;mem[13603] <= 30'b000000000000000000011001000000
                ;mem[13604] <= 30'b000000000000000000011001010000
                ;mem[13605] <= 30'b000000000000000000011001100000
                ;mem[13606] <= 30'b000000000000000000011001110000
                ;mem[13607] <= 30'b000000000000000000011111110000
                ;mem[13608] <= 30'b000000000000000000100000000000
                ;mem[13609] <= 30'b000000000000000000100000010000
                ;mem[13610] <= 30'b000000000000000000100000100000
                ;mem[13611] <= 30'b000000000000000000100000110000
                ;mem[13612] <= 30'b000000000000000000100001000000
                ;mem[13613] <= 30'b000000000000000000100110010000
                ;mem[13614] <= 30'b000000000000000000100110100000
                ;mem[13615] <= 30'b000000000000000000100110110000
                ;mem[13616] <= 30'b000000000000000000100111110000
                ;mem[13617] <= 30'b000000000000000000101000000000
                ;mem[13618] <= 30'b000000000000000000101101000000
                ;mem[13619] <= 30'b000000000000000000101101010000
                ;mem[13620] <= 30'b000000000000000000101101100000
                ;mem[13621] <= 30'b000000000000000000101111000000
                ;mem[13622] <= 30'b000000000000000000110100000000
                ;mem[13623] <= 30'b000000000000000000110100010000
                ;mem[13624] <= 30'b000000000000000000111010110000
                ;mem[13625] <= 30'b000000000000000000111011000000
                ;mem[13626] <= 30'b000000001000000000000001000000
                ;mem[13627] <= 30'b000000001000000000000001010000
                ;mem[13628] <= 30'b000000001000000000000001100000
                ;mem[13629] <= 30'b000000001000000000000011000000
                ;mem[13630] <= 30'b000000001000000000001000000000
                ;mem[13631] <= 30'b000000001000000000001000010000
                ;mem[13632] <= 30'b000000001000000000001110110000
                ;mem[13633] <= 30'b000000001000000000001111000000
                ;mem[13634] <= 30'b000000001000000000010101100000
                ;mem[13635] <= 30'b000000001000000000010101110000
                ;mem[13636] <= 30'b000000001000000000010110000000
                ;mem[13637] <= 30'b000000001000000000011100010000
                ;mem[13638] <= 30'b000000001000000000011100100000
                ;mem[13639] <= 30'b000000001000000000011100110000
                ;mem[13640] <= 30'b000000001000000000100011010000
                ;mem[13641] <= 30'b000000001000000000100011100000
                ;mem[13642] <= 30'b000000001000000000101010010000
                ;mem[13643] <= 30'b000000001000000000101010100000
                ;mem[13644] <= 30'b000000001000000000110001000000
                ;mem[13645] <= 30'b000000001000000000110001010000
                ;mem[13646] <= 30'b000000001000000000110001100000
                ;mem[13647] <= 30'b000000001000000000111000010000
                ;mem[13648] <= 30'b000000001000000000111000100000
                ;mem[13649] <= 30'b000000001000000000111111000000
                ;mem[13650] <= 30'b000000001000000000111111010000
                ;mem[13651] <= 30'b000000010000000000000101000000
                ;mem[13652] <= 30'b000000010000000000000101010000
                ;mem[13653] <= 30'b000000010000000000000101100000
                ;mem[13654] <= 30'b000000010000000000001100010000
                ;mem[13655] <= 30'b000000010000000000001100100000
                ;mem[13656] <= 30'b000000010000000000010011000000
                ;mem[13657] <= 30'b000000010000000000010011010000
                ;mem[13658] <= 30'b000000010000000000011010000000
                ;mem[13659] <= 30'b000000010000000000011010010000
                ;mem[13660] <= 30'b000000010000000000011010100000
                ;mem[13661] <= 30'b000000010000000000100001000000
                ;mem[13662] <= 30'b000000010000000000100001010000
                ;mem[13663] <= 30'b000000010000000000100001100000
                ;mem[13664] <= 30'b000000010000000000100010110000
                ;mem[13665] <= 30'b000000010000000000100011000000
                ;mem[13666] <= 30'b000000010000000000100011010000
                ;mem[13667] <= 30'b000000010000000000100011100000
                ;mem[13668] <= 30'b000000010000000000100011110000
                ;mem[13669] <= 30'b000000010000000000101000000000
                ;mem[13670] <= 30'b000000010000000000101000010000
                ;mem[13671] <= 30'b000000010000000000101000100000
                ;mem[13672] <= 30'b000000010000000000101001000000
                ;mem[13673] <= 30'b000000010000000000101001010000
                ;mem[13674] <= 30'b000000010000000000101001100000
                ;mem[13675] <= 30'b000000010000000000101001110000
                ;mem[13676] <= 30'b000000010000000000101010000000
                ;mem[13677] <= 30'b000000010000000000101010010000
                ;mem[13678] <= 30'b000000010000000000101010100000
                ;mem[13679] <= 30'b000000010000000000101010110000
                ;mem[13680] <= 30'b000000010000000000101011000000
                ;mem[13681] <= 30'b000000010000000000101111010000
                ;mem[13682] <= 30'b000000010000000000101111100000
                ;mem[13683] <= 30'b000000010000000000101111110000
                ;mem[13684] <= 30'b000000010000000000110000000000
                ;mem[13685] <= 30'b000000010000000000110000010000
                ;mem[13686] <= 30'b000000010000000000110001100000
                ;mem[13687] <= 30'b000000010000000000110001110000
                ;mem[13688] <= 30'b000000010000000000110010000000
                ;mem[13689] <= 30'b000000010000000000110110010000
                ;mem[13690] <= 30'b000000010000000000110110100000
                ;mem[13691] <= 30'b000000010000000000110110110000
                ;mem[13692] <= 30'b000000010000000000110111000000
                ;mem[13693] <= 30'b000000010000000000111000100000
                ;mem[13694] <= 30'b000000010000000000111000110000
                ;mem[13695] <= 30'b000000010000000000111001000000
                ;mem[13696] <= 30'b000000010000000000111101100000
                ;mem[13697] <= 30'b000000010000000000111101110000
                ;mem[13698] <= 30'b000000010000000000111110000000
                ;mem[13699] <= 30'b000000010000000000111110010000
                ;mem[13700] <= 30'b000000010000000000111110100000
                ;mem[13701] <= 30'b000000010000000000111110110000
                ;mem[13702] <= 30'b000000010000000000111111000000
                ;mem[13703] <= 30'b000000010000000000111111010000
                ;mem[13704] <= 30'b000000010000000000111111100000
                ;mem[13705] <= 30'b000000010000000000111111110000
                ;mem[13706] <= 30'b000000000000000001000011010000
                ;mem[13707] <= 30'b000000000000000001000011100000
                ;mem[13708] <= 30'b000000000000000001000011110000
                ;mem[13709] <= 30'b000000000000000001000100000000
                ;mem[13710] <= 30'b000000000000000001000100010000
                ;mem[13711] <= 30'b000000000000000001000101100000
                ;mem[13712] <= 30'b000000000000000001000101110000
                ;mem[13713] <= 30'b000000000000000001000110000000
                ;mem[13714] <= 30'b000000000000000001001010010000
                ;mem[13715] <= 30'b000000000000000001001010100000
                ;mem[13716] <= 30'b000000000000000001001010110000
                ;mem[13717] <= 30'b000000000000000001001011000000
                ;mem[13718] <= 30'b000000000000000001001100100000
                ;mem[13719] <= 30'b000000000000000001001100110000
                ;mem[13720] <= 30'b000000000000000001001101000000
                ;mem[13721] <= 30'b000000000000000001010001100000
                ;mem[13722] <= 30'b000000000000000001010001110000
                ;mem[13723] <= 30'b000000000000000001010010000000
                ;mem[13724] <= 30'b000000000000000001010010010000
                ;mem[13725] <= 30'b000000000000000001010010100000
                ;mem[13726] <= 30'b000000000000000001010010110000
                ;mem[13727] <= 30'b000000000000000001010011000000
                ;mem[13728] <= 30'b000000000000000001010011010000
                ;mem[13729] <= 30'b000000000000000001010011100000
                ;mem[13730] <= 30'b000000000000000001010011110000
                ;mem[13731] <= 30'b000000000000000001011001000000
                ;mem[13732] <= 30'b000000000000000001011001010000
                ;mem[13733] <= 30'b000000000000000001011001100000
                ;mem[13734] <= 30'b000000000000000001011001110000
                ;mem[13735] <= 30'b000000000000000001011010000000
                ;mem[13736] <= 30'b000000000000000001011010010000
                ;mem[13737] <= 30'b000000000000000000101101000000
                ;mem[13738] <= 30'b000000000000000000101101010000
                ;mem[13739] <= 30'b000000000000000000101101100000
                ;mem[13740] <= 30'b000000000000000000101101110000
                ;mem[13741] <= 30'b000000000000000000110011010000
                ;mem[13742] <= 30'b000000000000000000110011100000
                ;mem[13743] <= 30'b000000000000000000110011110000
                ;mem[13744] <= 30'b000000000000000000110100000000
                ;mem[13745] <= 30'b000000000000000000110100010000
                ;mem[13746] <= 30'b000000000000000000110100100000
                ;mem[13747] <= 30'b000000000000000000110100110000
                ;mem[13748] <= 30'b000000000000000000110101000000
                ;mem[13749] <= 30'b000000000000000000110101010000
                ;mem[13750] <= 30'b000000000000000000111010000000
                ;mem[13751] <= 30'b000000000000000000111010010000
                ;mem[13752] <= 30'b000000000000000000111010100000
                ;mem[13753] <= 30'b000000000000000000111010110000
                ;mem[13754] <= 30'b000000000000000000111011000000
                ;mem[13755] <= 30'b000000000000000000111011010000
                ;mem[13756] <= 30'b000000000000000000111011100000
                ;mem[13757] <= 30'b000000000000000000111011110000
                ;mem[13758] <= 30'b000000000000000000111100000000
                ;mem[13759] <= 30'b000000000000000000111100010000
                ;mem[13760] <= 30'b000000001000000000000001000000
                ;mem[13761] <= 30'b000000001000000000000001010000
                ;mem[13762] <= 30'b000000001000000000000001100000
                ;mem[13763] <= 30'b000000001000000000000001110000
                ;mem[13764] <= 30'b000000001000000000000111010000
                ;mem[13765] <= 30'b000000001000000000000111100000
                ;mem[13766] <= 30'b000000001000000000000111110000
                ;mem[13767] <= 30'b000000001000000000001000000000
                ;mem[13768] <= 30'b000000001000000000001000010000
                ;mem[13769] <= 30'b000000001000000000001000100000
                ;mem[13770] <= 30'b000000001000000000001000110000
                ;mem[13771] <= 30'b000000001000000000001001000000
                ;mem[13772] <= 30'b000000001000000000001001010000
                ;mem[13773] <= 30'b000000001000000000001110000000
                ;mem[13774] <= 30'b000000001000000000001110010000
                ;mem[13775] <= 30'b000000001000000000001110100000
                ;mem[13776] <= 30'b000000001000000000001110110000
                ;mem[13777] <= 30'b000000001000000000001111000000
                ;mem[13778] <= 30'b000000001000000000001111010000
                ;mem[13779] <= 30'b000000001000000000001111100000
                ;mem[13780] <= 30'b000000001000000000001111110000
                ;mem[13781] <= 30'b000000001000000000010000000000
                ;mem[13782] <= 30'b000000001000000000010000010000
                ;mem[13783] <= 30'b000000001000000000010101000000
                ;mem[13784] <= 30'b000000001000000000010101010000
                ;mem[13785] <= 30'b000000001000000000010101100000
                ;mem[13786] <= 30'b000000001000000000010101110000
                ;mem[13787] <= 30'b000000001000000000010110110000
                ;mem[13788] <= 30'b000000001000000000010111000000
                ;mem[13789] <= 30'b000000001000000000010111010000
                ;mem[13790] <= 30'b000000001000000000010111100000
                ;mem[13791] <= 30'b000000001000000000011011110000
                ;mem[13792] <= 30'b000000001000000000011100000000
                ;mem[13793] <= 30'b000000001000000000011100010000
                ;mem[13794] <= 30'b000000001000000000011100100000
                ;mem[13795] <= 30'b000000001000000000011110000000
                ;mem[13796] <= 30'b000000001000000000011110010000
                ;mem[13797] <= 30'b000000001000000000011110100000
                ;mem[13798] <= 30'b000000001000000000100010110000
                ;mem[13799] <= 30'b000000001000000000100011000000
                ;mem[13800] <= 30'b000000001000000000100011010000
                ;mem[13801] <= 30'b000000001000000000100101010000
                ;mem[13802] <= 30'b000000001000000000100101100000
                ;mem[13803] <= 30'b000000001000000000100101110000
                ;mem[13804] <= 30'b000000001000000000101001110000
                ;mem[13805] <= 30'b000000001000000000101010000000
                ;mem[13806] <= 30'b000000001000000000101100000000
                ;mem[13807] <= 30'b000000001000000000101100010000
                ;mem[13808] <= 30'b000000001000000000101100100000
                ;mem[13809] <= 30'b000000001000000000101100110000
                ;mem[13810] <= 30'b000000001000000000101101000000
                ;mem[13811] <= 30'b000000001000000000110000110000
                ;mem[13812] <= 30'b000000001000000000110001000000
                ;mem[13813] <= 30'b000000001000000000110010110000
                ;mem[13814] <= 30'b000000001000000000110011000000
                ;mem[13815] <= 30'b000000001000000000110011010000
                ;mem[13816] <= 30'b000000001000000000110011100000
                ;mem[13817] <= 30'b000000001000000000110011110000
                ;mem[13818] <= 30'b000000001000000000110100000000
                ;mem[13819] <= 30'b000000001000000000110111110000
                ;mem[13820] <= 30'b000000001000000000111000000000
                ;mem[13821] <= 30'b000000001000000000111001100000
                ;mem[13822] <= 30'b000000001000000000111001110000
                ;mem[13823] <= 30'b000000001000000000111010000000
                ;mem[13824] <= 30'b000000001000000000111010010000
                ;mem[13825] <= 30'b000000001000000000111010100000
                ;mem[13826] <= 30'b000000001000000000111010110000
                ;mem[13827] <= 30'b000000001000000000111011000000
                ;mem[13828] <= 30'b000000001000000000111110110000
                ;mem[13829] <= 30'b000000001000000000111111000000
                ;mem[13830] <= 30'b000000001000000000111111010000
                ;mem[13831] <= 30'b000000010000000000000000000000
                ;mem[13832] <= 30'b000000010000000000000000010000
                ;mem[13833] <= 30'b000000010000000000000000100000
                ;mem[13834] <= 30'b000000010000000000000000110000
                ;mem[13835] <= 30'b000000010000000000000001000000
                ;mem[13836] <= 30'b000000010000000000000100110000
                ;mem[13837] <= 30'b000000010000000000000101000000
                ;mem[13838] <= 30'b000000010000000000000110110000
                ;mem[13839] <= 30'b000000010000000000000111000000
                ;mem[13840] <= 30'b000000010000000000000111010000
                ;mem[13841] <= 30'b000000010000000000000111100000
                ;mem[13842] <= 30'b000000010000000000000111110000
                ;mem[13843] <= 30'b000000010000000000001000000000
                ;mem[13844] <= 30'b000000010000000000001011110000
                ;mem[13845] <= 30'b000000010000000000001100000000
                ;mem[13846] <= 30'b000000010000000000001101100000
                ;mem[13847] <= 30'b000000010000000000001101110000
                ;mem[13848] <= 30'b000000010000000000001110000000
                ;mem[13849] <= 30'b000000010000000000001110010000
                ;mem[13850] <= 30'b000000010000000000001110100000
                ;mem[13851] <= 30'b000000010000000000001110110000
                ;mem[13852] <= 30'b000000010000000000001111000000
                ;mem[13853] <= 30'b000000010000000000010010110000
                ;mem[13854] <= 30'b000000010000000000010011000000
                ;mem[13855] <= 30'b000000010000000000010011010000
                ;mem[13856] <= 30'b000000010000000000010100000000
                ;mem[13857] <= 30'b000000010000000000010100010000
                ;mem[13858] <= 30'b000000010000000000010100100000
                ;mem[13859] <= 30'b000000010000000000010100110000
                ;mem[13860] <= 30'b000000010000000000010101000000
                ;mem[13861] <= 30'b000000010000000000010101010000
                ;mem[13862] <= 30'b000000010000000000010101100000
                ;mem[13863] <= 30'b000000010000000000010101110000
                ;mem[13864] <= 30'b000000010000000000011001110000
                ;mem[13865] <= 30'b000000010000000000011010000000
                ;mem[13866] <= 30'b000000010000000000011010010000
                ;mem[13867] <= 30'b000000010000000000011010100000
                ;mem[13868] <= 30'b000000010000000000011010110000
                ;mem[13869] <= 30'b000000010000000000011011000000
                ;mem[13870] <= 30'b000000010000000000011011010000
                ;mem[13871] <= 30'b000000010000000000011011100000
                ;mem[13872] <= 30'b000000010000000000011011110000
                ;mem[13873] <= 30'b000000010000000000011100000000
                ;mem[13874] <= 30'b000000010000000000011100010000
                ;mem[13875] <= 30'b000000010000000000011100100000
                ;mem[13876] <= 30'b000000010000000000011100110000
                ;mem[13877] <= 30'b000000010000000000100001010000
                ;mem[13878] <= 30'b000000010000000000100001100000
                ;mem[13879] <= 30'b000000010000000000100001110000
                ;mem[13880] <= 30'b000000010000000000100010000000
                ;mem[13881] <= 30'b000000010000000000100010010000
                ;mem[13882] <= 30'b000000010000000000100010100000
                ;mem[13883] <= 30'b000000010000000000100011010000
                ;mem[13884] <= 30'b000000010000000000100011100000
                ;mem[13885] <= 30'b000000010000000000101010010000
                ;mem[13886] <= 30'b000000010000000000101010100000
                ;mem[13887] <= 30'b000000010000000000110001010000
                ;mem[13888] <= 30'b000000010000000000110001100000
                ;mem[13889] <= 30'b000000010000000000111000010000
                ;mem[13890] <= 30'b000000010000000000111111000000
                ;mem[13891] <= 30'b000000010000000000111111010000
                ;mem[13892] <= 30'b000000010000000000111111100000
                ;mem[13893] <= 30'b000000000000000001000101010000
                ;mem[13894] <= 30'b000000000000000001000101100000
                ;mem[13895] <= 30'b000000000000000001001100010000
                ;mem[13896] <= 30'b000000000000000001010011000000
                ;mem[13897] <= 30'b000000000000000001010011010000
                ;mem[13898] <= 30'b000000000000000001010011100000
                ;mem[13899] <= 30'b000000000000000001011010000000
                ;mem[13900] <= 30'b000000000000000001011010010000
                ;mem[13901] <= 30'b000000000000000001011010100000
                ;mem[13902] <= 30'b000000000000000001100001000000
                ;mem[13903] <= 30'b000000000000000001100001010000
                ;mem[13904] <= 30'b000000000000000001100001100000
                ;mem[13905] <= 30'b000000000000000001101000000000
                ;mem[13906] <= 30'b000000000000000001101000010000
                ;mem[13907] <= 30'b000000000000000001101000100000
                ;mem[13908] <= 30'b000000000000000001101111010000
                ;mem[13909] <= 30'b000000000000000001101111100000;

        end
        else begin
            state_reg       <= state_next;
            ptr_pic_reg     <= ptr_pic_next;
            num_line_reg    <= num_line_next;
            compute_out_reg <= compute_out_next;
            complete_reg    <= complete_next;
            spike_reg       <= spike_next;
            i_buff_empty_reg <= i_buff_empty_next;
            if (ren2in_buf) begin
                ptr_packet_reg  <= ptr_packet_next;
                packet_reg      <= packet_next;
            end
        end
    end

    always @(packet_out_valid, tick) begin
        if(tick) compute_out_next = {250{1'b0}};
        if(packet_out_valid) begin
            compute_out_next[249 - packet_out] = 1'b1;
        end
    end

    always @(*) begin
        ptr_pic_next    = ptr_pic_reg;
        ptr_packet_next = ptr_packet_reg;
        num_line_next   = num_line_reg;
        packet_next     = packet_reg;
        case (state_reg)
            IDLE:begin
                i_buff_empty_next = 1'b1;
                ptr_packet_next = 0;
                ptr_pic_next    = 0;
                if (start)
                    state_next = LOAD;
                else
                    state_next = IDLE;
            end
            LOAD:begin
                i_buff_empty_next = 1'b0;
                packet_next = mem[ptr_packet_reg];
                if (ren2in_buf)begin
                    ptr_packet_next = ptr_packet_reg + 1'b1;
                    num_line_next   = num_line_reg + 1'b1;
                end
                if (num_line_reg == num_pic[ptr_pic_reg])begin
                    state_next      = COMPUTE;
                    num_line_next   = 0;
                    ptr_pic_next    = ptr_pic_reg + 1'b1;
                end
                else
                    state_next = LOAD;
            end
            COMPUTE:begin
                i_buff_empty_next = 1'b1;
                if (tick) begin
                    state_next = LOAD;
                    if(ptr_pic_next > 2) spike_next = compute_out_reg;
                end
                if (ptr_pic_reg == NUM_PIC)begin
                    //complete    = 1'b1;
                    state_next  = WAIT_END;
                end
                else if (grid_state == 7)
                    state_next  = LOAD;
                else
                    state_next  = COMPUTE;
            end
            WAIT_END:begin
                i_buff_empty_next  = 1'b1;
                if (tick)begin
                    ptr_pic_next = ptr_pic_reg + 1'b1;
                    spike_next = compute_out_reg;
                end
                if (ptr_pic_reg == (NUM_PIC+4)) begin
                    complete_next   = 1'b1;
                    state_next      = IDLE;
                end
                else
                    state_next  = WAIT_END;
            end
        endcase
    end
    
    assign packet_in    = packet_reg;
    assign state        = state_reg;
    assign num_pack     = ptr_packet_reg;
    assign spike_out    = spike_reg;
    assign complete     = complete_reg;
    assign input_buffer_empty = i_buff_empty_reg;
    
endmodule