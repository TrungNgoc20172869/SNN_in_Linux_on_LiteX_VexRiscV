module neuron_grid_datapath_3x2 #(
    parameter CORE_NUMBER = 0
)(
    input [255:0] axon_spikes,
    input clk,
    input reset_n,
    input initial_axon_num,
    input inc_axon_num,
    input new_neuron,
    input process_spike,
    input update_potential,
    // output spike_out,
    
    output done_axon,

    output reg [29:0] packet_out,
    output reg spike_out_valid,

    input inc_neuron_num, init_neuron_num, shot, local_buffers_full,
    output nb_finish_spike
);
reg [367:0] neuron_parameter [0:255];
wire [1:0] neuron_instructions[0:255];

wire [255:0] spike;
reg [7:0] neuron_num_shot, axon_num;
assign nb_finish_spike = neuron_num_shot == 255;



always @(negedge clk, negedge reset_n) begin
    if(~reset_n) begin
        neuron_num_shot <= 0;
    end
    else begin
        if(init_neuron_num) neuron_num_shot <= 0;
        if(inc_neuron_num) neuron_num_shot <= neuron_num_shot + 1;
    end
end
// assign spike_out = shot & spike[neuron_num_shot];

// assign spike_out_valid = (~local_buffers_full) & shot & spike[neuron_num_shot];
// assign packet_out = (shot & spike[neuron_num_shot]) ? neuron_parameter[neuron_num_shot][29:0] : {30{1'b0}};
always @(negedge clk, negedge reset_n) begin
    if(~reset_n) begin
        packet_out <= 30'd0;
        spike_out_valid <= 0;
    end
    else begin
        packet_out <= (shot & spike[neuron_num_shot]) ? neuron_parameter[neuron_num_shot][29:0] : {30{1'b0}};
        spike_out_valid <= (~local_buffers_full) & shot & spike[neuron_num_shot];
    end
end

assign done_axon = (axon_num == 255);

always @(negedge clk, negedge reset_n) begin
    if(~reset_n) axon_num <= 8'd0;
    else if(initial_axon_num) axon_num <= 8'd0;
    else if(inc_axon_num) axon_num <= axon_num + 1'b1;
    else axon_num <= axon_num;
end








wire [8:0] potential_out [0:255];
genvar neuron_num;
for(neuron_num = 0; neuron_num < 256; neuron_num = neuron_num + 1) begin
    wire reg_en;
    assign reg_en = (neuron_parameter[neuron_num][112 + axon_num] & axon_spikes[axon_num]);
    neuron_block neuron_block(
        .clk(clk),
        .reset_n(reset_n),
        .leak(neuron_parameter[neuron_num][57:49]),
        .weights(neuron_parameter[neuron_num][93:58]),
        .positive_threshold(neuron_parameter[neuron_num][48:40]),
        .negative_threshold(neuron_parameter[neuron_num][39:31]),
        .reset_potential(neuron_parameter[neuron_num][102:94]),
        .current_potential(neuron_parameter[neuron_num][111:103]),
        .neuron_instruction(neuron_instructions[axon_num]),
        .reset_mode(neuron_parameter[neuron_num][30]),
        .new_neuron(new_neuron),
        .process_spike(process_spike),
        .reg_en(reg_en),
        .potential_out(potential_out[neuron_num]),
        .spike_out(spike[neuron_num])
    );
end

integer i;
///////Khởi tạo csram
generate
    if(CORE_NUMBER == 0) begin // x = 0, y = 0
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
            neuron_parameter[0] <= 368'b10101000101010101010011010001110101010101010001000001000111111101010010110100100100010100101000111001010010110101001110100000101110001100010000100010101010010001000001100101011110101000010011101110110000001011010100010101100111011011111100010001100010010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000000000000;
neuron_parameter[1] <= 368'b01011010101010101101010001010100110010101010101000000001110001011010101010001000011101011101101010101010000101011100001010101000000101010101001111011010100101010101011111101101010101010101010101110010101101010100010111010100101010101111010011010110001101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000000010000;
neuron_parameter[2] <= 368'b01001010001010010010010101110000100000100011101010100111010110100110010110101000110110010010111001010010101000100110011010111011011010101010000110101010101101011010101111010110101010110101101010000111011110101011101010101000000010110100101101111011110011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000000100000;
neuron_parameter[3] <= 368'b01001100110010010010010101010101010101101001001010010101010001010110100100101001010101010101001010010010100101000010101100010001001010010001101110110101010100100100000111000111010100010010010010111001001110010100010010001001101011011111011000000001001000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000000110000;
neuron_parameter[4] <= 368'b01001010011010101010101001110101110110101000101010101000010010101010011001011010110110101010010100001101010101011001101110100111011101010100100111011001010101010100011010010001010111011001010101011100000001010110101011010100111101011000101011100001101101000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000001000001000000;
neuron_parameter[5] <= 368'b00100100001000001010001010000110110110000000101100110101100101010000010010110101011001011011010101001010010101100111110101100001100101010100001101010010100010010111101000101010101010100101001010100101100010101010101010101001101110000001001110110000101111100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000001010000;
neuron_parameter[6] <= 368'b11010100000100010110101010111101101000000001111010101111011110101100101111001010101010000010101010101010101010101001111010101010101010101010110011001010101010101010101110110010101011101001101000100001110010101011011010111010101101011010111111110011010110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000001100000;
neuron_parameter[7] <= 368'b10110100101010101010000101001010111010101010100010110000101001101010101001011000000010100101001010000110010010101000001101000101010011010011000100110100001101010101011101010111010101010101011101110011001101010100010101010110010011110000110000011111101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000001110000;
neuron_parameter[8] <= 368'b01011010101110101010110110000001101010111101010110011100010011001001010101010101101100101001001111101011010101100011110100101010101001111100101110001010101010101010100000100000101010101010100010001111111010101010101010101001110011001111000001111001010101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000010000000;
neuron_parameter[9] <= 368'b00100111010101010110101011010010101001010000011010110101000000010100110011001101010101111010101010100001001000010011001010111100010100101001011100001010101011111010100000011110101010101001101010001111000110101010101000101000110011110111011010100001010011010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000010010000;
neuron_parameter[10] <= 368'b10101011000000110101101010111010001011010100010010101001101110101011011100101010010010100111100001101010101011011001001001100001101010010100110010110101010010101101011011111001010101010010010101011011100001010100100101010100010001001001111111010111010101100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000010100000;
neuron_parameter[11] <= 368'b10100101000110010100100101001010010110001001011010110100100111010010000101101001010101010100011001010110100101000100010110100101001100010100100001001001010010000101000011001000100101011011000110101100010110100010101010101110100100001000100011101010111011000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000001000010110000;
neuron_parameter[12] <= 368'b00100110010101010001101010101010101110101000101010100000001100101010101010101000010101010100101010101001010101010000101110101011110101010000010010011101101000010101011011110001010101111101010101111010110101010100010101010111101011111111010011011000110011110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000011000000;
neuron_parameter[13] <= 368'b10110000101010000100101000001010011010101001000010110000100101010010100110101011011001100011000000010110101001001000010101000101010010100111011001110100001101101011011001110111010000000100100101010110011001010100010101010111111110000100000100000100011000100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000011010000;
neuron_parameter[14] <= 368'b10111010010100110000101010101010101110110011110010101010110110101010010110101010101100010010111011101011010101011100101010101101011101011100011111001010100011010111100010010110101010111001100010000100110110101011101010101001100100011100010011111111001000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000011100000;
neuron_parameter[15] <= 368'b10100101010101000010100010100010010001010101000001010010101101010101010101010001001011110001010101010100001010101101011101110101011010101111101101100101011101101010100110011110100101100010101010100001110110101010001000101011100010011110110100100100101100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000011110000;
neuron_parameter[16] <= 368'b01111101010010111010010101010101100101001001101111010100010011100110110000110101010100001010001010001001000111010100010111001010111010101010010010001010101010101010101000010110101010101010101010101011101010101010101010101001111001011100100000111001110011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000100000000;
neuron_parameter[17] <= 368'b11101000101001011010100000010110001010100100101000000001100100101011000010100100000101010110100001001010110001010001100001010100101001010001001101110011011010110011010011111110011101101011011100011100011001010110100101010101000010010000000110000100010101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000100010000;
neuron_parameter[18] <= 368'b10101010100010101010101101010010100111101010011001000101100100000111011100010101000100100101010101010101010101010111101101010101010101010101011101110101010101010100011111011111010101010101010101011001011001010100110011010010011011000011000101000010111001010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000100100000;
neuron_parameter[19] <= 368'b01000110001110010010100101010100000110001010001010010100000000100000100100110101010101100101100101010001010101010001100010110101000101010101100011101001010100000111010011111001010100011101010110110011100111010100100011010101101001000001111000100101110100010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000100110000;
neuron_parameter[20] <= 368'b00111001010110101001010110100011100101010010100100101000001110100011011010111100110010000010111101101011110100011110111011110100101000011100110111001010111110101010101100000100101010101010100010100001111110101011101010101001111001010110001101101000101001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000101000000;
neuron_parameter[21] <= 368'b00110101010101101000000010110010010101010010100010001011000101000000001010001001011101110011010100101001100100010100010110110110100100010101101000001010000010100010100000010110101000000000101010100010100010101010101010101000101010110011001010111011001101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000101010000;
neuron_parameter[22] <= 368'b10101010001000101001011110011010100110101110010100101111011010111010001001010001101110100100100101110101001010111011011010110011010111101100001001001010001101010111110001000100001010110101000011100100011000101011111010100101010011110000111011100000010111100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000101100000;
neuron_parameter[23] <= 368'b01010000010001010010100100011101001000010101101010010100110001111100101010101010010111100011000010101010110101010011101100110010101000100011001111110111001010100101000001011001010100101011010101011111110001010100100101010110000100101000011100001111010011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000101110000;
neuron_parameter[24] <= 368'b10101011100001010101010101001010100001010101010101111010101110110101010100001111101010000011101101111011101010101010111011110110101000101010010011101000101011100010100000010010101010101010101000000111110010101010101000101010011001001100000010101110000000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000110000000;
neuron_parameter[25] <= 368'b10110101010101101010100000101111010101010101101101010010101001010101010110110000001001110110010101010110101110100011001111010101010100100101000011100101010101010110001010101010101101010100101010010000110110010101010100000001100100011111010100000111010110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000110010000;
neuron_parameter[26] <= 368'b01111000100001001010011010010111101010000000101001101001111000111101011010100100100000001111010101101010010011011110101001010010101101101011100111111100001010001100011010001010010100101101011111010100001000010100100011011010011010101010010000011011001001100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000110100000;
neuron_parameter[27] <= 368'b10110111001000101010010000001011000110001010000101001111000010011001000101010100011000101000110101010001011000100000010110011100010101110100110010010010101001010111100111000000001010110101000101101010000100101101011001010100010001001010110101001111010101100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000110110000;
neuron_parameter[28] <= 368'b10111011101010010010100101101010001000101001001011100011101111110010110110101001001110101110100001010010110101011000011010010000101011011100001010111100000010101111011111100011010111001011010101011001001001010110100011010101000101011000110000010000010110110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000111000000;
neuron_parameter[29] <= 368'b01000101010110010010100001010101111000010101101100010100000101010001000010010101000001111001010010101010100010100111110101001010101000101011101100000001001011101010101101110110111010101010101010100010001110111010100010101011100111110100000010010110001010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000111010000;
neuron_parameter[30] <= 368'b01111010101001011010010101010111001010010100101011100001111000101000000010100101010010111110000001001010010101011010101001010110101001001010010100101110001010110010011011111011010100101001010100011111101101010110100011000001011010101010111110001010000110010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001000111100000;
neuron_parameter[31] <= 368'b11010001010101010011001110101000011011111110101101001010101001011110101010110101101011111101100010101011100010101010110101001010011100101011011000010101001001001010010010111001010101010010011101110000100101010101000101010110101110000101101000010010100111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001000111110000;
neuron_parameter[32] <= 368'b01001011101010101011011101001101101010101010101000010110111110101010100111001010111010010001011111001010000111101001110101100100011101101010001011010101010010010101011101001101010101001011010101010011010101010100010011010100101110100011011101011010001001110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000001001000000000;
neuron_parameter[33] <= 368'b10110101000101010101001010101011110100010000100111101010001101010100101000010110101011111001101010101011101010101001010110101010101010101011101110001000111010101010101100111000101010101001101010100000110010101010101010111000000010110100000000111000010001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001000010000;
neuron_parameter[34] <= 368'b10111010001010010110110010101010100001101001001011000010100011100010110100101001010100010010001010010110110101011011110010101011010101011100100100101010101101010110001110001001110110110101010011001100011010101010101010101000011101000000111110111100000000100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001000100000;
neuron_parameter[35] <= 368'b11100100100000101010000100000110111000110010100001011100100001010000011011010000000000100001010100101001001000010100001100011010100110110001110011110101101000000101010010100111011000100101011101011110110101010100010001010111011110111100110000011111011000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001000110000;
neuron_parameter[36] <= 368'b10101000100100100100101111001010110100111010110010100001101101110100101101001010010010111001010101110100101011011010101001010001000010100101010000110101010000101010011100111111110101000010110000101010111010010100000010000101110100000001100000001111000100110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001001000000;
neuron_parameter[37] <= 368'b00001010101011010101000101010100000010101001010000100101000000101010101011000001010101100001101010101100000001010101101010101010100100010101100100011010101010110011010011011101001000100100011100000000111001110101010101010101010011000111100100111111110010010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001001010000;
neuron_parameter[38] <= 368'b10111010100000101001000101100011100110011010010100001111011110101111010101011010111101010100101110110101001011010001101010111010010110101100011010101010100101000111111000111001001010110100010001000101110001001011111010100110010110011011111001111010110101000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001001100000;
neuron_parameter[39] <= 368'b00110110101010010000110000010110010111101010101010111101111100010010101010010100001001101101101001010101000001101101110011010001010101010100101110000100100101010101010001111101000110100101010101110011110100110101110011010101110100011110001011110010011110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001001110000;
neuron_parameter[40] <= 368'b01011010101011001101010101111101101010101011010110000100010110101010101011100101010100010010101010101010001010010110110010001010101010101000100100001010101010101010100110011001101010101010101010000000010010101010101010101000001010101000100001100110100100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001010000000;
neuron_parameter[41] <= 368'b10100100101010101001001010001010010110101010001110100000101101010100010100100010001011000101010101001000111010101001100101010100001011000110001010110101010100001101011111101111010101010110010101011101000001010100110101010100111111101111100001010000100111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001010010000;
neuron_parameter[42] <= 368'b11111000101000101001001010101111110100000110100001101011101001110001001010010110100010100001001110101001011010111101101101101011010000101011011001110100001101011010101000010110110010100000111010011111010101011000010110101100111100010010100010000100010000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001010100000;
neuron_parameter[43] <= 368'b01001000010100001011010101011101110011000010101010010101010100000000011010100101010000101011010011001100010101111000000101011001010101010100101010000110100101010101010010001100001010101101010101110001110000101001101000110100111011001001101001010101010110000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000001001010110000;
neuron_parameter[44] <= 368'b11101011100110100100101101011011000101001011000010100001101000010110101101001011010010001011011010010100101011001010111001100101011010101101011100101000010000101010001100101111110101000010110010101100011111011100001010101011010010000101111100111101001110010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001011000000;
neuron_parameter[45] <= 368'b10111000000010100100101010111010110011001010010000100111000101010010101001000110010101111101001010100001011101010111111010101010100101010101111110101010100011010101010001010110011000010101010100001011000001010100010101010101100110001001011110010111101001000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001011010000;
neuron_parameter[46] <= 368'b01001010101001010010101010101000100111110101101010101010110110101010010101101010101000001010101011111101101001001001011010101001011101010000011100101010101011000101100100011010101010101001000011001011110010101011101010101011001001011010100111111011001010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001011100000;
neuron_parameter[47] <= 368'b00010010101010110101010010110010001010101010010100000010100110101010101010000000011001101010101010100100101001011011101010101010000000010101100100101010100101010101011111111111010100010101010101010011000001010101010101010110000110100011111110001101111000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001011110000;
neuron_parameter[48] <= 368'b11111001011100101101001011010100111100101010110000101001101011011010001001100010100010000111000010100101101010101011111100101011110110101001111011101010001101010010111110100110111011000000111010111111101101011000010010000111001111111110001110011100110111110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001100000000;
neuron_parameter[49] <= 368'b11000101101010101010001000101001110110101010101010101101000001010101010001000000100001100101010101010100010111101000100101010101011001010101100001010101010000010101011010100001010101010101010101111100000001010101110101010101011000110100101001010011110101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001100010000;
neuron_parameter[50] <= 368'b10011010010101111010101010101000101000010101001010101011111010101100110101001010101010000010101101011010101011101111101010101101010101001010101111001010110111010111111100111100100010101001011101010110100001100011101010101001101001010101110111110111000000100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001100100000;
neuron_parameter[51] <= 368'b00100010101001000010010100110010100110101010101101011111110000011010101000010000001101111100101000010101000000010001101010100101010101010101100100000101010101010101010111110001010101010101010101010011110101010101110001010100100110011111011111011110011110000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001100110000;
neuron_parameter[52] <= 368'b11000101011101011101011110101001111010110000011111000110011111011110101010101010111111101010101010101010101110111010010100101010101010101011001110001010111010101010101100011010101000101010101010000000011110101010101010101001010010000110101111100110001101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001101000000;
neuron_parameter[53] <= 368'b10110101000000010100101010101010010101100001010100011010101111010010000101010101010010110101100010110100000010101111000101001011011100000010010101000100101011101010101001101010100001101010101010000110000010101001100100101000110110010001001010110000010011110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001101010000;
neuron_parameter[54] <= 368'b11011101010101001001001000110100101101010010101100100101011011010101001010010010110101001011011010101001011011000100010101101010100100101001001000001010101011011010000000111110111010100000101010000000101110111000101010101010001011101100111100011001001110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001101100000;
neuron_parameter[55] <= 368'b00110010100000101011010100110010000110001010010100001001100000101010110101000101001001111110101001010000010001010000101010010101010001010101101010001101010101001101010111001101010101010100010101111110001101010101110101010111100111111000011101011100100111010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001101110000;
neuron_parameter[56] <= 368'b10101011010101110100101011101001000101010000000010100011101110100101110101011010101010110000111100110101011001001111001010101011010101001110110101001010101011100101101110000010101010111011100001101110111010101011001010101000110011110010101011100111011001100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001110000000;
neuron_parameter[57] <= 368'b10110111010101000101101110101010000101010100010100001011101100001100101001010110001001100000001000100101001000101110001010111101010110000110100110100010100101010101101011010001101001010100101001100010100100101001111100000110101000000000010101110011111111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001110010000;
neuron_parameter[58] <= 368'b00101010101010010100101010101011100110101001000010101010010010101010111000000000010100001000101010100100010100000001011010101010100100001100110010001010101010000111100110000110101010101001100010000001100010101011001010101000100000010100101110111100111110010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001110100000;
neuron_parameter[59] <= 368'b01010100101000011001011001100100010010110100110101100010010011011010100101010110110101110010101010101001010010000010110010001010100101100111000100001010101010010011100011110100101011111101101010000100010010101011011010001010000101000010000011110111110111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001110110000;
neuron_parameter[60] <= 368'b11011101001100100100101101100100110101001010110010110100011111010101101001011010110010000001001010100100101101001110010001101010110010101010100010001100101101101010101110011110111010100101101010000000100010101010001010101011001010011011110000111000111101110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001111000000;
neuron_parameter[61] <= 368'b10110101010100101001001010111011010101010010010101101010101001010101000100010010101011011111010101001000101010101010101101010101100110101001100101110101010101001010101110001010010101010100101010010000111101010100010100000111111000000001011110010100101101110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001111010000;
neuron_parameter[62] <= 368'b10111010101010010000100001101011000110101101101000001011101010100010110110010011001010111110101001010101010100101111001010000101010101010110000001111100100101010101011011000001010111010101010101110011011101010101010101010111010110010010001000000111101101000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000001001111100000;
neuron_parameter[63] <= 368'b10100011010011011001001010101010000100100101000101101010111010001010010010010100001010000110101101001001010010101010001110010100100101100010101111010100101011010101101000011101000100101001001000000100010001101001111101010000100001011011111011101001010010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000001001111110000;
neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
    else if (CORE_NUMBER == 1) begin //x = 1, y = 0
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
                neuron_parameter[0] <= 368'b10101010110101101010010101001000101011111010101000000010101010101110100010101010101010101010010010101010101010101010110111011100101010101000000100010100010100001100010100110011010010010101010101010101001011011001000110001001010101000111100101001011001111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010000000000;
neuron_parameter[1] <= 368'b10101011011011101010000001101010101001000000101010101000101010000111110010100000010011000001010011001010000101010101010111000101000100010101010111010101010101101101000100011100100101010100101000000110011010011110001000101010111101100110111100110100111001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010000010000;
neuron_parameter[2] <= 368'b10010011101110110110100101000010010110111110010101111001011001101010110010001001000101011010101111001010001110110100101010101101101010101001011110101001110110001010101101010010101001010001000010010000011010111101010000001001000010101010110101110010100101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010000100000;
neuron_parameter[3] <= 368'b11010101010011001011010110101011101100010000101001001010101010011101011010110100001010101010100110101101010100101010101000000010100101010010100001000100001010100101010000100000010010101001010101101000100011010010101001010100111000100100101110001100010000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010000110000;
neuron_parameter[4] <= 368'b00101010111100110101010010001010100011011001010101000010000101011100101101010101010101010101010010110101010101010101010101111011010101010101010101010011101100000000010101010100001010101000101000010101111010101010001000000010101010101010101010001000000010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010001000000;
neuron_parameter[5] <= 368'b01010110111111001001001001010000101011110100100000100101001010101100000010101110000010101010110100101010101110101010101011011100101010110010100111001001011010101010010111000101101100101010000001010001010011111001110100010100010101100101010101000101101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010001010000;
neuron_parameter[6] <= 368'b00010101100000101001010101000101010100101000010101010101010101010001001001110001010101010111100100101000010101111101001010111010101100101010101010101011101010101000101011101110011110001010100010101011110101101000101100011111111010000001101010111001001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010001100000;
neuron_parameter[7] <= 368'b11000101011001010101011000101101010111010101010100100100010101010101010100010010101101010100000000010011010010100101010101100101010101001010010101010011010111010100001101010101011101001011001100110101010101111100101010010101000101010100011110100000010101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010001110000;
neuron_parameter[8] <= 368'b11011010000000101010001011110101000010101110100010000001010100101000101010110101010101011010111110101011010101010100101000101010100101010100101010100100101010100100000010101000000110001010100010100000101101101010101010101000001010010001101010101010101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010010000000;
neuron_parameter[9] <= 368'b11010100001111010101010110101100000010110111010101001011010001111100111101000110101000001100000110100101001010111101000000010010110001001011100100011101101000010110100011101011011110000000010010100010101101100010110101011000001000100111101010101100001010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010010010000;
neuron_parameter[10] <= 368'b00101010010001001010101010101010101011010111101000001010101010101101110010100010101000010010000111001000100010010101000001001100100000010101010101000001010000000100010101000101010010010101000001010101011000001101100101001000110011100101111110001000101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010010100000;
neuron_parameter[11] <= 368'b00100100110011011001100001010010011010010010110000101101000011111010110100110010010010101010111011010101100101001011001100100101010101010100100000110001010101010101011011000001010101100101010100101000000101010000001000010010101010010000000100000101001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010010110000;
neuron_parameter[12] <= 368'b01010100011111010101010101010101010101011101010101100001010101111000000101000101110101010010101010101010001111110000001011011010101000101010101010101011011000101010101010101010100010000000101010101010001010011101101010101110100001001011011000101010101100000000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010011000000;
neuron_parameter[13] <= 368'b10101010101000101001011010100010101010011010100101001100010110111001001010110110101001011010101100101010101010000101101010101110101010101001010110101011001010101010010101010010101100101011100101000100001010111110101001010101100010101011111010010101011010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010011010000;
neuron_parameter[14] <= 368'b10101010101000101010101000101011010100111010101001110111010101010000111101110110110101010101101011010000010001010101010100101001000100101101010101110010110111010110110101101010101101111010001001001011101010100001000110100101001110101011100010011010010100110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010011100000;
neuron_parameter[15] <= 368'b10001010100101010100100001000010001000010101000010010100000000101101110110101001011000001010000010101010100101000111001001010110101011010000011000010101001010101001000000101101000010101010110101000100000100101010101010000000100001000101101010101010100000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010011110000;
neuron_parameter[16] <= 368'b01101011110010111010100101010010110111011010101011010111011010010011101010101101010101011000010111001010010101010111100111010100101001010111111100100000010001101001001100010000000001011010101100111110001000011101101100010100100010000111010100000110101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010100000000;
neuron_parameter[17] <= 368'b01010101001001010101010101010101010101100101010100010100011000101001000100000011001010100010000100101010101100001010101000101110101010000010101010101001001010101011001010101000101110101010100000001010010100111100110000000101101001011100011010100110000000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010100010000;
neuron_parameter[18] <= 368'b00000010010111100000001001001010101011000001000011101100101010101111110010001001001010101010000110100111010010101010101001011100100110001010101010100111011011001011000110010001010010100100000001010101001101011010000110100101010101010100101010010110001101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010100100000;
neuron_parameter[19] <= 368'b01000101101001001010110010010101010100110010110100101101010101010011011101000100100101010101101101010101000110100101010010101001010111101010010001101111100100011000001011001010101100010001101100101011011010100101011011110110101010101010010101001101001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010100110000;
neuron_parameter[20] <= 368'b01000010101000110101111101010100010010111101010000100001010011101010110101000001100101101010101110010110001010011011100110111111010010101010100110011011111101010010101010110100100011110111011010110101010101100000111011001101000110011001000111110100110010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010101000000;
neuron_parameter[21] <= 368'b00000101100101111001101011010000011011000000110100101001011010101111100010010010101010101010101011001101100010101010101011110010110011011010101010101111001011100000001010100000110111101101001101100100000001110010110100010101000001000100101011000101010101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010101010000;
neuron_parameter[22] <= 368'b11010110101110101000101001010100010010111110101001101001010101101010010010101010100101010100101101010010101010010101100010110011111010101011001010001010101100011011101000011110101011010101110100100110010010110001010001000010100100001010110101010010001110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010101100000;
neuron_parameter[23] <= 368'b01000111001101101010010110101001011110110010110000001010110101011010000101010100101011010110101111010001100110101100001010101101010011001010010100101111010100011100101101000010101101010101111010110101101010110100110110011101010110001110110010101001110101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010101110000;
neuron_parameter[24] <= 368'b10010110110010110001100111010001001000101101101011100101010110100110110110100000010100001010101011010111011001010010100111110101010001110101101010100011100101010101010110101100000011100100010111001010011111000001010000010110101000010001000001011000001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010110000000;
neuron_parameter[25] <= 368'b10101011101110110001000000010010010100100111010101000010010101010101011100010101010101010101010000010101010101010101010100010011010001010101010101010000101100111010100101010100011010101010101010111001011100101000000000100000101010001010101010101100000010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010110010000;
neuron_parameter[26] <= 368'b01000101010010110101000010010000101111011100010011000010101000011101101011000101101001010100000111111100010110010100010011011101010100010101001110011100010101010101010110101001110010010101010010111010101111011001011110101010000000000111111101101010100100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001010110100000;
neuron_parameter[27] <= 368'b00010101010111001101100111010000010100010101101011011011010011101010110010100101101100101010101010101011010110101010101010101010101101011010101010001011001011010100101000100001001110100111010010000000110100101010010101001000010101000000101001100110101010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010110110000;
neuron_parameter[28] <= 368'b10010100110110010101101010101101010011011101011000001010010101000100001101001001101101010010010100101001011010110100101001011010110100001001001010100101001010010100100100101010110110101001001010010001101010000010101000101001010000101010101010110010110001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010111000000;
neuron_parameter[29] <= 368'b00010100101101010000110001001011010011010101010001010110101101011100110101010001001010110101000100010101010110101101011111011010110101001010010101001000010001010000101001010100001111110000001111000101001001000010100101010000110101101111001000010100000001010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001010111010000;
neuron_parameter[30] <= 368'b10101000110110100101001000101000100101011001010110000010101011010111111100010001010010101001000111010101010101010110010101000101010101010100101001010100010101000101111000010100100011110111011011011101011010010010001001000101010101010001101000010101010001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010111100000;
neuron_parameter[31] <= 368'b10110000101011101001001000011010001011100110100001100001100100001111110100000010100010010101010011010100101011010101010101010101010110001001010101011100110101010100100101010100011101110100011110010101010010110001001001000010010010101010101001010010101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001010111110000;
neuron_parameter[32] <= 368'b11001010011001110100101010101010101011000001101000101010101010101100101011000000101010100010100010000100000001010000000001010100010101010101010001001111001011000101010100100100000010111111110001010101101010010010101101100011010001110110101001101001110001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011000000000;
neuron_parameter[33] <= 368'b10010010011011100101000010010101101001100001010010101101000000010110011000001010010101000100011101101010101001010100110101101110101010010100001001000000001010101001010010101101000110101010001000001010101111001000101000001010000001000000101010101110000001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011000010000;
neuron_parameter[34] <= 368'b10101001101000110111011010101000010111001010100010101010101101001100001010101101101010010110010100101010001010100001010111011010101010101011010100011100001010101010101101010000000010101011001001110100100011001110111101010011010100101111110101010101010011010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011000100000;
neuron_parameter[35] <= 368'b00100101000101111000010101001000011000000011000101010100101010101011110101010100111010101011001001010010000000101010111101110100001010101010101001110100011011101010101000010001110111000010000011001010100011001100010001010101010110000000110101010101010000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011000110000;
neuron_parameter[36] <= 368'b01010011011110100001001010010001101001101010100010101101010000000010101010100010010100000011111110011010101101010000100111111101001010110100000010101011010100001001010000000101111000110010100100000100010010011101001010010100000100101011101110001100100101010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011001000000;
neuron_parameter[37] <= 368'b01000000011010011100101000110101010010101101010001000010010101000101100110101000101101010110000001001010100110110100111011001101100010001001010110101101010100001010100100010010111001011100001011010101101011101111100000101001010101001000110110101010101101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011001010000;
neuron_parameter[38] <= 368'b10001000010110101010001010001001100000101010101000101100101110111011110111100000010010101011101101010000010101001010101110100101010001010100101010111001110101010001000010101011101001010000000011001010101110111101010000000010101010111010111100010110101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011001100000;
neuron_parameter[39] <= 368'b00001010010101101010101101011001001000000011101001010101100010100010101101010101011010101001101000110101010101101010110100100010010101011010100101010000011001010101101001000010010101100100000010100100001001000010101101001001100010111001000001111010001010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011001110000;
neuron_parameter[40] <= 368'b01000001001110001000000010110101000111001100010110101011010101010010011101101010101001010100000101010100001110100101010001010101010111010010110100101101111100010101101010010100001010010011001100101001010101111001101010101011110011000101111010100010101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011010000000;
neuron_parameter[41] <= 368'b01101010101011100110110000000110101011000011010001000010001000101100011101010010101000010100010100010101010000100101010101001011010101110011010101000100001001111011011101011100000110100011101101111101101010000010000011110000100100101111001000101110010010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011010010000;
neuron_parameter[42] <= 368'b01010101001100010100100101000010111100100101010101001110001100101010110101010001001010110101101110010101010100010101010000011010010101010101010101011011101001010101010101010101001010101000110000010100111000110010101000101000100100111111101010101010101010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011010100000;
neuron_parameter[43] <= 368'b00010001101011101001010011110001000100110010110101001000000001111010101011000100101011101010101010101101010010101010101010100010110101011010001110000111001011000101101011100010001110101101010110100000010110100010000001011100111000100001101010010101101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011010110000;
neuron_parameter[44] <= 368'b11110000110000110001001001011000101000100000101000100101100000101000100100100000010110101010111011010100101011011010101101100100010110100101101010110001101001010101010100001001000001100101010101010100001100001011010100100010000100010001101010010100100101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011000000;
neuron_parameter[45] <= 368'b11110100000001000101000101001010001100110111010001001100100000010011101101011101010010100000101010101111100101001010101000101010101010110101101011100010001010101011010110100010101110100000000000010010001110110011101100000101001001100000001111010101010000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011010000;
neuron_parameter[46] <= 368'b10010101001110010110000111000101010100010001010100111001010101010001110101000000100101010101001010110100001100100101010010101011111101101010010101101011101010111010101001001100001110001000110100100110011010110000110010111110110010101110101001101010100000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011100000;
neuron_parameter[47] <= 368'b10101000111000101010101010101010101011010010100010100010100000100100011000100000101001010101010001010100110010010101011001010101010101101101010101000101110101010001010101111110010101110110011101010011100100010001000101010001000100100010100101010001000101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011011110000;
neuron_parameter[48] <= 368'b10101001110110111110101110101010101000101010100001010101001010110011101000000001010100101011101001010000110101010110101010110101001110110101001010101000100101000010000010111010101000010000001010100000110000111100000100010011111010010010111000111111010001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011100000000;
neuron_parameter[49] <= 368'b00011000101010101011000100000001101010111110101011110010101010111001111010101000010000101011111101101010101000010110101110100000101010101001011010111001110100001010100100101011101001010101000110000010111110101101010111010110101010101011010101000100001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011100010000;
neuron_parameter[50] <= 368'b01000001010000100101000110101001010111011100010010010010010101011100001011010010101101010100110110101101111010010101000001011010100000010101000011000101001010111001010010100111010010101010101001101011101111011010001010101000001011010101101010101010100000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011100100000;
neuron_parameter[51] <= 368'b00001010111111010100101010101110101011010101101010101010101010101100110110101010101010101010110111100110101010100001011011010101000100000000010101000101010001010001010101100000010111000101010101010100001011010110010100000100010101001111010110000000101001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011100110000;
neuron_parameter[52] <= 368'b01010110001111101101110010100100010001011010010101001001000011011101000001010010100000010101111011010101101011010001010111100101010110101100010101011010110101001010010100000000011001010110101001000100001011000111010010110101011010101111010101010010110001010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011101000000;
neuron_parameter[53] <= 368'b00101010001111001010110000100010101101010010101011010010100000110101101010100101001010000111010110101011010100101111010001010010101001010010010101001100001010101101010101010100110110101010100001000101110010001011001010001000110011100101001010101001101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011101010000;
neuron_parameter[54] <= 368'b01011001001000010101001101000101100110110101010010010101101000011010110100101001010010100001001001010010100101010101010100111101011010101101010101011010110100001010010101010101001001010000001001010101000100101101001110100101000101101011010101000010101010100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011101100000;
neuron_parameter[55] <= 368'b00111010010111000001000001011110101001010101100111010011001010110110110010010010100100101000111110100101000001010010101111111110010000010101001011000001001001100110010101101010010010100001001001010010101111010011100011000101001000110101000111010001010010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011101110000;
neuron_parameter[56] <= 368'b10101101010100101000010100101101010100111110101101000011010101010101101001000000110101010101001011110000010101010101011110100000010110010101000010111011100101010101000000110010001010010001110110101010011000000001000101001111001010010011101001011000101110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011110000000;
neuron_parameter[57] <= 368'b00100010110111110101000100000001011011100111010100001010000010101101001111001010010010001010010100100110101101001100100101001100101010010100101110110001011010101001010001010001111011101010100001100001101111001100101010000010000000010000001010101100100011000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000000000000001011110010000;
neuron_parameter[58] <= 368'b01010111101001011011010100000100011010001000101001000001101000101010001010101010101010101110111110101010101010101010111010101010101010101010100010101111001010101010110011101010100100101010000100100010001011011001110101010101000011111110000101010101011110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011110100000;
neuron_parameter[59] <= 368'b10101001110011000011101101001000001100110111010011010100110101010110001100101100010010010101011000101011001101001011010110101110001010110101100101011010011010100110010011010101001111101101010101011011010101110001110100000100101101010000000101010111010010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011110110000;
neuron_parameter[60] <= 368'b10100100110010110101101001000101010010101011010010101101000001001011000101101010010101000101101101010110101001010001100110100101010010100101000010101011110101001010010010001010111101010100101011000100011011111101011011000111000100011011110101110110110101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011111000000;
neuron_parameter[61] <= 368'b00101010111101000101010100001010101001000011000010010010101010110101011100110100001010101001010100101010100010100000010101011110101010101011000101011000011010101010100101010001111110101010101001011000101111011110101010010100010101101110110110010101010101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000000000000001011111010000;
neuron_parameter[62] <= 368'b01011001000110101010101010010100011000111000101010100101011001011011101010101011010101000100101111000010100101010010111010101101101010010101001110101011010010001101001101000010111100011000100010100101100010101001100100001100000100001011111110100101100011010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011111100000;
neuron_parameter[63] <= 368'b00001001001010001011000011010010010100100111010100100101010101010001001101011010110101010101001101010101001100010101010110101101010010101011010100011010110101011010101100001010101001010110000010000010001000100101011010010010100100101011010101010000101010100000000000000000000000000011111111110000000011111111110000000010000000000000000000000000000000000001011111110000;
neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
    else if (CORE_NUMBER == 2) begin //x = 2, y = 0
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
            neuron_parameter[0] <= 368'b01011110100011001000001101110101001010001010111100110101010101101011100110000101010100110110101111010100110100010101001010101101000001001100101000101010101101100010101010000011101010111100101010101001010100101011110101101010010101010101101011111110100101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100000000000;
neuron_parameter[1] <= 368'b10100000010101011100110110001100001010100001010011001010001100101010101011000101110010101010101010101100001100001010000110101010110000110010101001010110101011101110101010010101010100101100101111000101010100010100001011100101000001011000000110000101010100100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100000010000;
neuron_parameter[2] <= 368'b01010101010101010111011101010101000110010101011000010101010100001100000101011101010101001110100001010111110010010110100011010101010111011101101011010000010101010101111110100101000101011101011101001010010011010101001000110100101011010000110110110101010010100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100000100000;
neuron_parameter[3] <= 368'b01010010101010011011110001100001101010101111110010111001010100110000010001101011001101011010000000011010000100101100101010001100101100100011010010100011101010111111000101001010010101010011010101010000101011110001010111011101010010110111010101010000000011000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100000110000;
neuron_parameter[4] <= 368'b10111110101011011011000010111000101010000001001110100110101010100101101100001000111010001011010110101101001010101010011101000000111110100111100000110101000011011010110101010101010100100000100001010100010100101001001100110101010101011010100010111011010101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100001000000;
neuron_parameter[5] <= 368'b01010101010111010110111101000000000101011100100110011101000000000101000010101001010000000010100001001011000010100010101010101001101011100000001010101010001110000111000010001010100000001111011101010010101011011000011000111101010110100100000101111010101001010000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001100001010000;
neuron_parameter[6] <= 368'b00100010110100101010001000101111011011011000100110101111111001100011110111111010011010110110101111001011001110001010011010011100101010101000101001101101010110011010100010100110110100101010101101100010010011010100110011010101001000110111010101101111010100100000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001100001100000;
neuron_parameter[7] <= 368'b01010100101101010100100000010101001010000011000110100100010100101010000101101000101001010010101100011001100000100100101010110101101100101000011010001101000110111001100101101010010101011101010101010110010000001101000000111101010010001000010101010011000101000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100001110000;
neuron_parameter[8] <= 368'b10000001010010001010101010101010100001001100100010111001000000000101000101001011100010001010100101000000101000001100101010100101100100100001000010101010011111011010010111001010101101001100101001010101001010010100110010101000010101010101010111110010100101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100010000000;
neuron_parameter[9] <= 368'b00000000101000100100001101010101010010101110011000000100010101001010101001110110100101010110101010100111001010000000011010101010110100101100100101101010101001011010101010000110000011100101101010001100111011010000110110001001010101000101010111000010101100100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100010010000;
neuron_parameter[10] <= 368'b10110010101010101010100010001010010110000100001000000000101001010101010110001011001010010101010101001000100110101001000101010100000101001010100100110101010100010100101010011000001100010010100011100101001101000101001110000110110101110001010100101101101001010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100010100000;
neuron_parameter[11] <= 368'b10010100101010101010101010000101000001000001010010111001010111010101000000111010100011011001010101111110101001100101001001010010110010100101011010101001010100111100010100101010101100010010010101011010101010110001010011110100110010101000010111011011010001100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100010110000;
neuron_parameter[12] <= 368'b10100001010011101010110110100110000101000110100011000011100010010100101010100101000011001001010010101000010100010010100101001010111011010001100111010100101011110101100010100100001010101111010100101100110100101011010100011011111110000010101101011111110111100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100011000000;
neuron_parameter[13] <= 368'b10001010100101010110001010010000100000000101011001100100101011010101010101010111010110101101011001010100110110101010010101010100010001010010101101010001001101110100001010010101110110101100010010101100010101001010101000101010111001011010100011100100101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100011010000;
neuron_parameter[14] <= 368'b01011100010101011010000001011101101001000101001000000100001010110101110100010000001010101001010101000100111010101010100100010100010010001010101000010101011101101000101010110100110110001100001010101111000010101111001111101011010101001010110100101101110101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100011100000;
neuron_parameter[15] <= 368'b00011101001010111010001011010000010100101000101010100000010111010010101111001110000101010101001010010101101000010100010010101000111100101000010100011010100001101010100100001100101001101100101010000100001011100000110011001001000000000010100111000000101001010000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001100011110000;
neuron_parameter[16] <= 368'b11011010100101001010101010100110001011010111011110101010010100101011010001010010101101010110101011000111101010000000101010101001010110101010011000001010101111001010101010011101101010111101001010101001110111001010101110101010100101010010101100101100101000010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100100000000;
neuron_parameter[17] <= 368'b01100010010100011011010100000000100001011000110110010011101010000100011011111000100110100100010100101001000110101010010011010100000100001011101001001001110110001001000010100010101101010011010101011011001010110101000100110100101111101011010101010011010010110000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100100010000;
neuron_parameter[18] <= 368'b10101011100010101011001010101010101000101010101010101010101010000100101010101010101010010110000110101000001010101101011011001100110010101010010100100101101110111010101101010010010110110110100010110101111001011010010011001001000101010100101011111010101111010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100100100000;
neuron_parameter[19] <= 368'b01001010000010111010110100001000101010001110111001001010001010010010000000100100101010101101011000010000010010101000110101000100000001011010101011010101010000100110101010011001010101010010111010001001000001010111001101101011011010101001010100111100001100110000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100100110000;
neuron_parameter[20] <= 368'b00101000101010101000010000010000001010100010111101100100000010101000000011111100000111010101010100101010000101000111010101010110111101010010001001010101011010101100110100000101010101000110000000100000001001010101010010010001010000101000110101100001010101000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100101000000;
neuron_parameter[21] <= 368'b10010011001010001110100001001100100000000110000010010001110100101001010001001010100110100010101011000101001000000011001010101011101010110100010100101010101100001111010101001010101010110101000000010101010101101010010010101001010100010101000011000100100101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100101010000;
neuron_parameter[22] <= 368'b01010101000110101011111101111100100101000000111010110111010101010101101110110011011001010001010101011011111110100101101011010101001010010010101011100000010110101001101010101011100101011010000110101011101000000010111100000010101011110000111010101001000000000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100101100000;
neuron_parameter[23] <= 368'b10101010101010101010101010100010101010101001001101100011001010100101010101010010100100101101010101000100101000010010010101010100010100101010111101001001010001011000001101010100000101101001100011000101010101010100101000010100110101011001000010000011010101010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100101110000;
neuron_parameter[24] <= 368'b01111001101010010111110111000110011100001010011101010100100000010101101011100101011010010101010100101010010101000110100101010100011001010100000100010101010100110101010000100010110101010010110101010001101010010101010101010101010010101010010101100101010100100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100110000000;
neuron_parameter[25] <= 368'b00010001010101110110111100000100010001010101000011011101000101001000010101000101010100010010101001010111110101010100001010100101001001010101000100101011010100010111010010101010100101001110111100101000101011010000110011011010100010100101101011011100100010100000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001100110010000;
neuron_parameter[26] <= 368'b00010101101010111100000010010101010010101001100011001000110001000111101100100101101010000011010100011011110110101010101101011000011111001010101010110100100101110000100010111001011010000001110100001000000010100010001001001010011111001001001100101100101101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100110100000;
neuron_parameter[27] <= 368'b10101000101010101011001010100010000010101000111010101000101100101100100010101010101101010010001010001111101000010101101110111010110110110001010100100000011111111001010101010110010101011100000101010101010101000101110011010001010101010100000001010011001101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100110110000;
neuron_parameter[28] <= 368'b10001010101011011001100111110000101010000101001010000100001010101101010100000111010010001001010101010100101100101010000100010001010010100010110001010101010001101010101000010101011110110001101010110100010100001001001011101011010101001010101100110010111101010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001100111000000;
neuron_parameter[29] <= 368'b10010001011011011001111100000100010101000110100110011101000001101011001010110001010110100110101000111011100110011011001010101101101101011010101000101001010100010001000011111010100100001111010101010010101011010100110011010101100010101101010101010111010011100000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001100111010000;
neuron_parameter[30] <= 368'b10101010101010101010100100101010101010101010111100011110001010101010101001110101001010000000101010111010110010101000010101001101010001000001010001010101010001000111001010110001010101010001111111101001010101010101001111001010101010000001101010101000000110100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100111100000;
neuron_parameter[31] <= 368'b11000001010101010101110000101000110001010100000001011000100001101000000100010101010001010010101010010110110101010100001010101001001101010101010000101010100101110101010101010010101011000101010100110001001010100010110000010110000010100000100011101001001101000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001100111110000;
neuron_parameter[32] <= 368'b00001110101010111000110000010111100000100011101011001000010010110101011011101111101101000001010101001001000110100001100101010110100111001010100111010101011010101100101010001101010100110011101010101010110101010101001011001111001001010101110100101010110001100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101000000000;
neuron_parameter[33] <= 368'b10101010100001110100001010101000100010110110010100101010100010010011000011010110100001010001000011011001010100010101000010110001111101001001010100101001000110100100010101010110100010000010010101010100101000000001111001010101010100100010000011010011000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101000010000;
neuron_parameter[34] <= 368'b10101101000101001010001000100110100010110100001010010100001010101101000101001011010000111010110101010100101011010000101001010101010000110001010010110101010111001010100000000001010101010001000110011101010101000111101111001000110101010110000010101010001001010000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001101000100000;
neuron_parameter[35] <= 368'b10101010010100110100010100000110101001001001001101010100000010110101000100010101001001101011010100011001110100100010100101010010011101010100100011010101101000100101001010000101000010100011110100101110100101101010110000110110001001000010101011110111010100000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101000110000;
neuron_parameter[36] <= 368'b00011101101101110110111101010101011110011011011101110101111010010010100101000111010100010101100100010100011101010101010100010001010101010101010001010010100101000011001010000101101011110100010110101010001110110011101111001010101011000110111000101100101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101001000000;
neuron_parameter[37] <= 368'b01010101000110110100000100000111001100101011011001010101010100110010100001110100000101010101001000010110100000010111110110101011011000110101011101010010101101011110110100110101101001110101101000100011011010100101000101111010010001100000100110010000101010010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101001010000;
neuron_parameter[38] <= 368'b10001000101010101011001010100010010010101011101110101000001101101010101010111010011100010100100100101010001101010101010101010100100110110110010101010101010011110010011101010101010101001001101010110101000101011010001100111010010100010010101010111111001010100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101001100000;
neuron_parameter[39] <= 368'b10000011101010001011000010100000100110101010100010100010010001110010101010101010101010100011010110101011001110101001101111010010101110101010100110110101111010001010101111011011010101001001001011001110100101010101101110100101111100100101010100010111010010110000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101001110000;
neuron_parameter[40] <= 368'b00011010101010100110010110010010010110100010011100000101000001010100000011001000100101010101010101010011010011110101010101010101111001000001010100100101010110110101010101001010000101010110011101000000101000000101110000011010101010101000101011100011101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101010000000;
neuron_parameter[41] <= 368'b01000100001100010100101010010000010101010001000010100101100011010000000000000010111000101101001010000101101000101110110110100001010100100010101001011000100101011010010100100100001010111100101010011000010010101010110000101010001101001010101011000110101111010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101010010000;
neuron_parameter[42] <= 368'b10010011101010000101011010100010101100100010101111101010001001011010110010000101101010010100101111101000110011110101011001000101101101000001010101101111010110100100110101010010001011000011111101010101101000000001110001010101010010100000011101101101010101100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101010100000;
neuron_parameter[43] <= 368'b10101010101010101001110010010100001010101011001001100000010000010010001100101100001111001101010101001000110101010001010101010100010101010000000111010101010010111101110000010101010100001011110110010101010100100000101101010100101001001010101010001011010010010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101010110000;
neuron_parameter[44] <= 368'b00101101000100000111001010001010100001011101001000100100001010101010000000001010010000001010101010000001001000001000001010101010000110100100110110101010101011011010010000000001101010101101001001011000010100101010101011101101000101010101001010111100101000110000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101011000000;
neuron_parameter[45] <= 368'b10001001010100010000011001000110101010100001010001001101010010111010010101101001100101001011010101010101100101010110000101010001011001010101010000010101011001100101010101001001010001001000110001010111000100000101101110101000110010011010100110010001001111000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101011010000;
neuron_parameter[46] <= 368'b01000010101101100100000100001000000010100011111001010110000000010110101111010101100110110101011010001011110011100001010100100010111011010100100101011010010000000100110000010100101100110011100110010001011010000100011101010101010010101001101011001101010100100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101011100000;
neuron_parameter[47] <= 368'b00010000101010101010000110101000000010101010101100010010000000001010101010101100101001000100101010101010101010100100011010101010101010101110100100001110011010111010110111000010100111000011000001010101011011100101010100110101000101101111010101010010000101010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101011110000;
neuron_parameter[48] <= 368'b10100001001010101001110010101000100101001010111100101001101010010100101010011010101010101101010010101010100000100000110101101000111000100011100001010010101011111000011010110101001010101100000101010010010010101010110100110101011101001000000001001101010110100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101100000000;
neuron_parameter[49] <= 368'b10010100010010100100001110101100010101000000100110111010110101010000010101011110101010000101100100000011101010101101010010101111000000101010000000101010001100111010101010001010101000000110101010100000101010111000010010101010100010100000000001001100101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101100010000;
neuron_parameter[50] <= 368'b00011010111000011000100111011001101010000011001110000111011101001010110110000100110100010110101001010100111001110101010010110101010011000101010001101010101101101110010101000110110101010100001001000100011011010011011111011000000101000000010111011010101001010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101100100000;
neuron_parameter[51] <= 368'b01000100001001100110010100110110011100110100011001000011010101010010001010100100101101000101010010001000010010100100000101010111011101001010010100010110100110110111101001010101010011001010011010101101110101101011101001101010101011010010101010101100101100100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101100110000;
neuron_parameter[52] <= 368'b01001000101010100000010110101100000100100010111011100010110001011010101011110100100001010100101011001111010111000101010010101011111101010101010101101011011000010101010100000110101010100110010101000010101011000000010001010100100000100000010111011111011010100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101101000000;
neuron_parameter[53] <= 368'b00000000000101001000000101000110001101010101001001100101001000000101010110010110101010100101010100001001010010000001010100010100010101001010100101010000010000000110100001010100101011110010011010100101010010100001101001101010000101001010100010011110101000010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101101010000;
neuron_parameter[54] <= 368'b00001100000010101010011010011111010101010100101011011101000011010101011100101001001001010001010101010011110001010100101001010101001011010101010010101001010100010101000100101010101011011010111010001001100010101111011000011010010110101010101001111010101000010000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001101101100000;
neuron_parameter[55] <= 368'b00000101010101110110100100000000000101010100010110011011000000000000010001111010110000011010101001010110101001101000001010101101011010101101010010101010110101011011011100001010001011011100001111010010100101101101001101111100101011010011010100100101010010000000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101101110000;
neuron_parameter[56] <= 368'b00010001101010111010001011100110000110101010100110101100110100110010101000111011011000010001010100101000001000010100000101000101101010110001010010010111010100010101010110101001010101010011011111001010101001010101001010000010100010101001011110101001111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101110000000;
neuron_parameter[57] <= 368'b01010101100101000110010001010100010101010001101101001000000000000100001011010100101110100001010010110010011010111010010101001010001101001010101101011010101000110110101010101100101010101010010010110010101010101010110100010000001010101101101111000101101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101110010000;
neuron_parameter[58] <= 368'b10000011101000011111111001011010001010010101110001000101101001101001100111100101010101000110100010011010110111010101011011010110110111010101010101100101010010110101010101001011010100010110011101000000101001011001111100001010101010100010101011101110101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101110100000;
neuron_parameter[59] <= 368'b01000001010001101000100101010100000010010101010101010101110000001010010000000101110100001000101010000111110010101010100010101010011101010010101011011010101011111110101010100100011010101100000010101001010101110010101100101010010101010100000010101110101100010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101110110000;
neuron_parameter[60] <= 368'b01000000000000011011101000010100100000110011100110101001111010010110010000011010100101101011001100000110001001000110101010011000101010100001011010101001010111111010010101001010100100011101001101010100101011100101001110100000010100100100010100101010001010010000000000000000000000000011111111110000000011111111111111111110000000000000000000111111111000000001101111000000;
neuron_parameter[61] <= 368'b01010000000000101010110101000001010101010011111011010101001010001001001010010100011010100000110000101001010010101010110110001010110001001010101100101100001110110100101010111000100110111010010010101010010010101010000010101010100101000110101011101010101001010000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101111010000;
neuron_parameter[62] <= 368'b11000001000101010110011010110010100011010011100101011011111010100101001110011010101010101010010110101011110101101010101101000101001001010100101010110101000110100101001010101011010100011011110101001000101100000100110000010110011010010101111010001101010101000000000000000000000000000011111111110000000011111111110000000010000000000000000000111111111000000001101111100000;
neuron_parameter[63] <= 368'b01010100101011110100010101010101010100100011000011100110000100010110101100011000101001010001011010110011010101000010100101101001010101010010101011010110100101100001001010101101101000001010110100101000010110101110000100110110000010101001110110010101011000100000000000000000000000000011111111110000000011111111110000000000000000000000000000111111111000000001101111110000;
neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
    else if (CORE_NUMBER == 3) begin //x = 1, y = 1
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
            neuron_parameter[0] <= 368'b01011001110001111100110010110101000101010101010010010010100101010100010101011011100011110100000011100110001111000010100100101101001010101110001011000100000010101010010010100101110100101010101011111011100100000010101010101011001011000101001010100000000011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000000000;
neuron_parameter[1] <= 368'b10000101000111000101010000110111010101010101010101100111101101010101010100010101001000100001010101000001010101111101010101010100010100010111000101010001010010011010011100011001001000101010101001001001100100101000101010101100000000010000110010100010101001010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110000010000;
neuron_parameter[2] <= 368'b11110110101010101010101001010000101010101010101010101100010110111101101010101010001100011101011001111010101010001100010101010101101110101011100101010100110001111010100000110101100010010101101010000101010010101000010110101010100000101010100000001010100010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000100000;
neuron_parameter[3] <= 368'b00001010101110001100100110010101111010101010101101101110011010101010100010010101000110101010100001010001010101001101101001010001010101000100011010100101100001010100010101101011011000110100001101001110100100101001010010111001011011011000101101101000001010110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110000110000;
neuron_parameter[4] <= 368'b11011010101010101010101001110111111010101010101010101101000110101010101010101010101010011010101010101010111011110001011010101010101011010100000101101010101111101101010111110100101000000111010101111111010000010110011101000110011101001101011010111101011101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001000000;
neuron_parameter[5] <= 368'b00111110011011100111001000111100010101010101010010011000000101010100000101000101011110110001000000000101010101001011010110010000010001010101000101001001101001000100010001011001001100101010101101001000110100011010101010100101100010001100101010101010100011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001010000;
neuron_parameter[6] <= 368'b11111010011000110111001110111000111001110101010000111111101101011001010110001110101011010110110100101010101111010101010110001010101010100011011110110100101010101111010011000010001010100010001101001111001010001000010010001100010100101010010001000101001101010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000000110001100000;
neuron_parameter[7] <= 368'b00011010100111000101010100000011110101010101010100100100000001010100010101010101110010101010000000100101010100001011101010100000010101010101101010100001010110010101011100001011000110101111010111110010000100110110100101011000101001010001101010010101110100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001110000;
neuron_parameter[8] <= 368'b11100101110101001100111110110011001110010011100110000100111011011101010110101011010001001010100001001010101000000100101010010111101010101001110110101001000010101010101001011010100110001010101010101001101010000100101011011110101010101000110010100110111000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010000000;
neuron_parameter[9] <= 368'b11001110010101010101001100111100110101010101010100011100100101010101010101010101001011100011010101010101010101000001011100000001010101010101000100100100001001010101010110010010011000101001100101010000010000000010101010100100000010000000101010101010010110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010010000;
neuron_parameter[10] <= 368'b11101101010101110100100101010110000101010111110111010010101010001100001010101001001000001010010000101010100010100010101011010110101001011000101000101100010010100101100000110010100100101011110001010011001010000110100101000110010101001001001010110111001001010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110010100000;
neuron_parameter[11] <= 368'b10011101010101010101110010011111010011111101110101010110001001001010100100010101101100100100101010000001010000100101001010101001010100101000110100001010110101001010101000111101101010000000101010101011010110101001001010001000000100001010100000101001001001100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110010110000;
neuron_parameter[12] <= 368'b01101010101010101010101111001000101010101010101010101001011110101010101010101010101010011100101010101010100111000100011010101010010101010111011010110010101101000101010101000010000101000110000101001111101111010111101101011110011001001101010010010011010111110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011000000;
neuron_parameter[13] <= 368'b00111111111010101010001010001110100101001010111011001001100000010101000011101100110010100001010100100100011111110001010101010010100010010101101101110101011110100001011000010100010101001010010101011001000001010100111001010011010100101101010000100101000110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011010000;
neuron_parameter[14] <= 368'b01100100101000110010001000011100001000101010101010011101001101101010101010101010110111010110001010101010001011111100010010101010101011101010000110101010101011001101011111010011010100100010100001100101000001010100010010100111011001010111010101010000001001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011100000;
neuron_parameter[15] <= 368'b10101011110111001100110110111001101010101010101010100111010010100100101000110101101010101010000001101010001100110110101010010100001011101100101010100101010010101010100111101010010101001010101010111010100101011100100000101011101110010100010010001000101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110011110000;
neuron_parameter[16] <= 368'b10100001100101001100110100010000010010000001000110101011010110001110000100111011011000011010100000010111000110001010101010000101010001001100001010100010101001000101001000101010101010100101000101000010100010101010011001101101010101000110101101011110110100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100000000;
neuron_parameter[17] <= 368'b00001100011001010101001100001000010101010101010101011000001101010101011000011010011010100101010000101001001000010101010110011101010100101001100101011100011001011010001010010100100000000000100010100001010010101010101010101101000100101010101010101010111010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100010000;
neuron_parameter[18] <= 368'b10010011101010101000110110100001101000101010101010101010111111111100101010101010111111111111010000111010101011000000000101010101010110001010100100000111010101010110101011101101010101010101010110100000001010011001010101011100100100101000101010101010110000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110100100000;
neuron_parameter[19] <= 368'b01000010110101100111000011101110111011010100110101110001001100100010100001010001010001101010101000110001010101000110101010100010000001010110011010101011010010100001011110101010110101001011000101000000101001010100100001011000101110101000010111000100000010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110100110000;
neuron_parameter[20] <= 368'b01110010101000100010110110101101110101010101001010101010101100010101010110101010011011111000010101010001001101111010101100110101100010011000101010001110010110001010110110101010100001001011111011100010011010100100100101001111101011110000011001110100111110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110101000000;
neuron_parameter[21] <= 368'b01011100010111010111001100110110010101010101010101010001110001010101001001010010010011100101011100100110101010001100010100010001101110101001000101011001100110101010101010110110100001010100101010101000011011101001011010111010101000100000100101101010101110010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110101010000;
neuron_parameter[22] <= 368'b10101011100111001000110110000001110000101010101010101111000110101010101010101010110110101010101000011010101010101100101010110110101010111010011010101110010110101010100111101010100101010100101010011110111011001101011010101100101010011100100101001010111110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110101100000;
neuron_parameter[23] <= 368'b01111110110101010111001101001100010001010101010101010101110000010110100101010101100101101011000010100001010100001011101010101010001101010100001010101000100010000100110010101010100101001011010001000000101011010100010100101000101010101001101101010010000010000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110101110000;
neuron_parameter[24] <= 368'b01110100010001100101110011000001010111011101110111010000000101001010100101010101001001100100101010010101010100000111010110101001001101110110011101001010100000010101010010010100101011011000101001101001010010101100000010100111000010101010110010101011111110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110000000;
neuron_parameter[25] <= 368'b01111100010111010101011110000001010101010101100110011000000011000101010100101011010001100111010100001010101000011110110101010100101011101011100001010101001010101100100000110101010100001010110111101001010100000100100001010011101100001010010010010110101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110010000;
neuron_parameter[26] <= 368'b10000111011010110011001011001010000101011101010010011000110100010101101001000110110110110101010110000101011101101001010101011001000001010010101100110101000110100110010100111100110100101010010111101000011011010010101010010110001100100101101001101101010111100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110100000;
neuron_parameter[27] <= 368'b01110001110111010101011011011011110101010101010101001101101101011001010101010101011100100010101101010100000101101111101011110001010010110100011010101010100100010000100010101010100010000011100101011010101011000101110010100100001010101100100010101010010110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110110110000;
neuron_parameter[28] <= 368'b00101101000010111000100111100001001000101010110111000111010010011100101010001101000110000110101010101101101010010110101001101010101001001010101000011010101011001000101001110000010010101101000010101111010101010010010100011110011001010101101011100111101101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111000000;
neuron_parameter[29] <= 368'b11000010101110001010111010011100101010101010101100100110110010101010101010101010011011001010110100101010101010110110100101010111101010000011111011110101010000001110000101101101011100010110001010111110010110011101010111001011111101000101100101010100001101010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000110111010000;
neuron_parameter[30] <= 368'b01000000010101011100110110110001010001101100010010000010011101011110101000001011010101110110101010110111000000011101001110101000000001011000011100011010101000010000101000110001001010011000001011110001101110101001000010101011000110111010100000001010100110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111100000;
neuron_parameter[31] <= 368'b00000100101010101010101001100011111010101010110101001010001101111010100011100100010101110000010011000001011101011010010101011101010101010111011010100000010001010100001010100000101001000101000101100010101010001010101011100101101010101000101010101110010110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111110000;
neuron_parameter[32] <= 368'b00010110101010111010101101011111101010101010101011000011000010101010101010011010110100001110011010110001011011010010110101101000110100000110010001010010101011010101011000010101011010001011010101010011101101001100101101110001010001000100111010010100100101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111000000000;
neuron_parameter[33] <= 368'b00001110011010110111001000000100000111011101001100111011110100010100010110101010101000100101010100001010101011000011010101010010100110100110101101010101100000011010000100010000000010100001010101101000000110101010010110010011000000101010110101000101000000000000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111000010000;
neuron_parameter[34] <= 368'b01111001010101010101110101000110101011010101000100111111010010001010010100011010110111000010101000001001101000000101001010101100000010101001010000101000010011101010100101011010101011010010101010100100101110100111001010101011001010110010010100101010101010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111000100000;
neuron_parameter[35] <= 368'b01101101110101010101010000001111001111010101000100110000000010101010010000110101001000101110101000010010110100111101101010100101101001011000110101101010010000110101101000110010101001001011010100110001001010110100100010000101100000101010010010001010111010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111000110000;
neuron_parameter[36] <= 368'b00110011101010101000100010000010111110101011001001100111100110111110100111010101111001011001011111101001010111110000000101100110110101010100001011010110001001010101011000101101011100010101010101001110100101000001010100100110101010001110100101101001000110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001000000;
neuron_parameter[37] <= 368'b11010010101111000100110101001111110101010001011101100001011101110101010100000010000010111011010101010010011011011001000001010001010100010011000110010101010101010100001010010001010101000101011101011000000000010010101001001100100100100000101010101000110110110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111001010000;
neuron_parameter[38] <= 368'b00000001110101011100110111110011001111010010100100100100100010101011010001001010111100101110101101000110101010000111101010100101011010101011011100101010010000101010101010111010101000011010101010011101001110110101101010011010100110100011010110110000100010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111001100000;
neuron_parameter[39] <= 368'b00001010101110001010110101111110101010101010101010100110110110101010101010101010100010101010110100000010101011010110100101010110101010111110001010011001000110101010100010101111100100010000101011101010100000100001010000000010101010001010110101001100001110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001110000;
neuron_parameter[40] <= 368'b10110011010101001000110011110011101000101010100101110011110010101111111010101001000001101010011100101011001000101110100101010010101010011001001010001100100010100011101110101010100101001001000010100011110101010100100100101010101110000111011010010010100110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010000000;
neuron_parameter[41] <= 368'b11011100000101010110001111000011010101010101011101001010010001010110000101100100000111000111110010010010011010011011011010101001001100101010000110101010101001010100101000011010001010100101011010011101010001001010110101101001010101000100101011010110101101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010010000;
neuron_parameter[42] <= 368'b01011101100010101010101110111011001010101010110110100000001010101010101111001110110000001110101010110100111010000001110010101011110010001000110100010000101011011101100000010101100010101101001010011111010101000010110101101011110101000101101011010110101001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010100000;
neuron_parameter[43] <= 368'b11010010101111000000111100100010111010101001111010101011000100101010000101101010000101111001111001010110110011000001010001110101011000001001100111001000110101111110110110100101111011010010001110111000010100100101101001011000000101010000010111010100110110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010110000;
neuron_parameter[44] <= 368'b10100010101010101010101001101001101010101010101010100100001111101010101111011110110100011110101010101000010101000100011110101001000101000101010111010110101010001101010101010101010110001010100101010111010101010110100011000111110001011101010010101001100101110000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000000111011000000;
neuron_parameter[45] <= 368'b10100110011011010101010110001100010101010101011101111010010100010101010101010101000100100001010101000101010101111011000001010100101000010110100111000001000010101001011110101000010100101000100101001011010101001000000110101001101101010100101110101010101010110000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111011010000;
neuron_parameter[46] <= 368'b00010011100011001010110000111001101010101010100001100111100010101010111111111000110111001010101011101010101111010100100011101010101101000110011010010000101010110101010110100101000010101001001101010011101101011010101101000101010011010101001000001101100101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011100000;
neuron_parameter[47] <= 368'b01011100101110001010101101011011101011101010100111000111110010101100101010101010000100001101010000101010101010000100110100101010101000100001000101011010101010111001100110010101000101011000110011101101010101010110101011010110010101010001010010000011111101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011110000;
neuron_parameter[48] <= 368'b10001010101001100010111111010011101010100000011010100100001110101010110110110011110010011000101011101001010111001001010100101010010101010101100101010101001011010111011110010101010010100101100101010100010110101011010111100011111101010000000101011011001101010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000000111100000000;
neuron_parameter[49] <= 368'b00011101011101110111001100010111010101010101010101011010011001010101100001010101000001100010000010101101010100000110010010101010001011011011010000100100101110101010011110001011001010100110101010111101010000001101000010110011100101100000010101010001000101010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000000111100010000;
neuron_parameter[50] <= 368'b10010001010101110101010100001000000101010101001000111011010011010011010010110001000100101001101111001011010100101011101010101010101101001100101010101010000010000101110101001010101101101110110111011100101000001100011010101000101010000100001111101010100110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100100000;
neuron_parameter[51] <= 368'b10011101010111010101110011101111000101010100110101010110011001010101011010101101011010000101010000101010110000100101000000010110101001101011100101000000011010100000101010011000000000101010110010111001101000000010100101000011100101000001001001010101011001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100110000;
neuron_parameter[52] <= 368'b01011100010001010111010011000110010101010101010101111000001100010101001010011101000110100101000100101001010100010101011011011010100101011010110000110100101000001001001100111001011010101100100011111001010100101010010011001010100101100010101101010010100011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101000000;
neuron_parameter[53] <= 368'b11100110111000110011001010110111000111101001100000010110101001010010100110111010111111010101101010101010101011110000010010101010101010100010000111101010101010001010010001010100000010100000001100100001010101010100010111000010011011010011010101010100011001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101010000;
neuron_parameter[54] <= 368'b00000010011010100010110110011010110100011011000110100001110101110110100101010100000111110011011011010101011101011010100001110101000010010110101010000100000010100011010010101000010100101001100101101010110101001010100110101001101001010100101000101010101110100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111101100000;
neuron_parameter[55] <= 368'b10111101010101010101010101000011000001011010110101010101011001010100101001010101011010100101011010101101011010111111100101001010010001101000111110010100101101000000101010011001000110110100000010111101101001011011011001101110110010100000100100000010011100100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111101110000;
neuron_parameter[56] <= 368'b01011010101010101010110100011110111010101010011110100100011110101010100111111110010100011010100001010100011011001001111100010101010101011110000001010111001001010100101110100100110010101001010100110010011010101010100101010101000101111010101011010101011010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111110000000;
neuron_parameter[57] <= 368'b11110100011011110111001101110110010101010101010101011111101101010010110101010101010001100101101011000101010101111111010110100101011001010101000011100010000000000101010001000110001000001010101101010000100111001100101010100100101010001000101010101010110101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111110010000;
neuron_parameter[58] <= 368'b11001010100110001000110100010111101010101010101010101100110110101010001000101011010011001100101101010100100010001000101010111101010010001000011010001010101101000110101100101010101010100000110010001010101010100011011111011001001110001110001101011100100110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111110100000;
neuron_parameter[59] <= 368'b11001101011010110011001111101101100101111001101101011010001001010011101010101110111111010100001010101010101110101101011010101010101011100000110101010000101010100100011001011000000010101000100101110101001001001010000111100100010000010011100101011000011001010000000000000000000000000011111111110000000011111111110000000010000000000000000000000000001000000000111110110000;
neuron_parameter[60] <= 368'b10111101010101011010110011101001000000101010010010011100111010010010101001000011111010100101011010100101001010000100000101101010000011101001111000010100101001001010101111101010011010111100101010010000101001001011001010010111100010001110100100101001001101100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111111000000;
neuron_parameter[61] <= 368'b11100001010111011100110100100000100100000010111101000010111000010011001010100101001111001011000000101011000000111100100001010010100101101001110010100101011010010101101010011010010100100101010100001000101000010010010000101000110010101000101000000010111000010000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111111010000;
neuron_parameter[62] <= 368'b01111101010101110101110111100001010101010101010101011111010101010101010101010101001101110011000101010101010100000111101000000101110101001100001000100101010110111010111110110010001000111011110011101001010001101001011010101011101100101000101101101011100010100000000000000000000000000011111111110000000011111111111111111110000000000000000000000000001000000000111111100000;
neuron_parameter[63] <= 368'b11010101110111010101010001001000110101001001001110010110111011000101011100101010000100100101011100001010101000011110100101000000101010101000100101001000101010101010100100111001000000010010110010110011010000000101101011100011101111010001010110100010011010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111111110000;
neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
    else if (CORE_NUMBER == 4) begin //x = 0, y = 1
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
neuron_parameter[0] <= 368'b01101000101010101010100001000110011001101100110000101000101000100111111111101011000001110000110110001111011111001011011001000010001001111001010001000001100011100001000001010010010010001000001000010001110111110000011110001001010110110001101010100000010011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000000000000;
neuron_parameter[1] <= 368'b10110110001100011110111001101101100100001100000110100111111001000010001010101011100000001010000110010011001100100101001010111000101010001000101110110110011000001110001110001100001100111100000000100000011011101111101010010011100011101000010110001000100000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000000010000;
neuron_parameter[2] <= 368'b01000010010000110101001100011001100001001000110001001101001001010100110111110010110001111010000100001101011101001000011010001010100000101001011001000101100001101001100000000000001111000010001000100001000000000100001101000011101000001100011110010100000110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000000100000;
neuron_parameter[3] <= 368'b10111010001010100010101110101010011010101011101011101000101000101010111010101010101010100011101000101000101010111010100000001010111011001010101010100010101010111010110010101011001110101010101011101011100010101110101010101010101010101001101011101000101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000000110000;
neuron_parameter[4] <= 368'b00011011000101100101111001111000010111000010101001010101000010011011111010001010000110100010110011100000000001111010001000110000101010011000111010100011101111101010000001110000001100011001001001111110100000101101111000011110010111010000010000000000100001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000001000000;
neuron_parameter[5] <= 368'b10100001111100101000000010000000011000111011010010001000010011110010000000100000000110100010001001001000100000110000100001101101010111111111000011101011110101100000111000100011110010101100110110011010110110011010000010100001000011010010101000000010010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000001010000;
neuron_parameter[6] <= 368'b10111000000010001010000001000110100001100100001010101000101000100101110000101001110000110000001110110110110010110001000000010010011101001011100100001010110100001011101111100001000110111100101000001010100010010001100010110010010111000000000000001110101000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000001100000;
neuron_parameter[7] <= 368'b01010000011100001000100000010100011001011000100100000101000000011001111001111100001010100010100000001001100011100010000101000011100010101000011001100001100011010111010001100010110011001010000110000010100101010001000000011001010011100010100000001100011101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000001110000;
neuron_parameter[8] <= 368'b10101011111011111010110100010001000111100010110010001000101100100101001000001011110000100110001010110110011100111100111011111101101000011110000101101111011000010100010011100010001000001011100010100010101000001010001001100010010010001000011010100111000110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000010000000;
neuron_parameter[9] <= 368'b00111000001101011010101111100110111000010000000000100101011010000000001000001010011100000111101111111110000001100000000010111001000001100000100100000000111000100010100101100010010010001000110100101110110111101110100010001100100010100001101011010100111010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000010010000;
neuron_parameter[10] <= 368'b00100101100010101010001011101111001010100001011011111000111100100010111001111000101011100110101000000110110011000010100000111010111011011000100000010000101110100111010110010010000000011110101011101101111011101111101010001000110111110000100011010100110011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000010100000;
neuron_parameter[11] <= 368'b01100001001100011110011001100101000000000100000100100111111001000100010010111001010000001011001010011011001100000111000010111100111000001000101010010110011000001110001110001000001000101100000010001000111010101001111010110010111011101001100010001010100000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000010110000;
neuron_parameter[12] <= 368'b10000011000000010111110010011001000010100010100110101110011101100100110001000011100001001010001110111111011100001001101010101100001000100011001010010010001000000000001101011100000101000000110101001101000000000110000000101100101000001001001011110000010011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000011000000;
neuron_parameter[13] <= 368'b11101100110010111001101000111000001010110111011000010000010100001011001100101100101110011001111001100000110010110010000100001101111001000010111110010010000000001110001110011101100000100000000110101100101011000100001101001110100000101001011010100001101101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000011010000;
neuron_parameter[14] <= 368'b00010100000000000110100101110010010100011000000011110000100000101010111110011010100001111001000101101001001010100010010010100000101000101110101000001110100010101011010000101010000110011011011011010001010110010001110011010100101010111100110000001100001000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000011100000;
neuron_parameter[15] <= 368'b10101110110000010000001000001000010000001011010000000000110101011010000000001000001010000001011001001001010100000110110100000100010101111101000100101000110101110010111000100001110011101010110111010011110110001011010010111001000100000010001000010000010110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000011110000;
neuron_parameter[16] <= 368'b00101010110110100001101000001000101011000010100001001000011011001011110111011101110000110101000010110011000111101100010010111010010101001111000011001010010111001011101000110000100110111100111001011010111010010001010010110110010111000010010010001100000100010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000100000000;
neuron_parameter[17] <= 368'b00010001111000001000000101000110010001001100110000100101000000000011100000111001001010011010100000001001000110100000000011000010001110011001111100101001100010010111110110101011111011011011100010011010111010111111011010110011010111100010000011001100011101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000100010000;
neuron_parameter[18] <= 368'b00101110101010100000000100011010100000101101010010001010101011000110010010010001111001000110100110100111110110100001111010101011101000011110101100110101001110100100100111010011111000001011111001100011000001100011100110000010010110111110001000000100101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000100100000;
neuron_parameter[19] <= 368'b00010010000101001010110011100101011000011000000011000111101010011001101100100110011101000000110011110110001011010010010110110000110000110100100101001100001011110100100000101010010010001111000000000000000101000010101111001000101000111010101001110101111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000100110000;
neuron_parameter[20] <= 368'b00100110100011101100010000011011100001100100011101001010101100100111101101101010100011110010101110000111111111001011001000100010111000101001101010100000100110111010100110010010000010101011101000011100001001100111111110001010011110110011101100101000011011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000101000000;
neuron_parameter[21] <= 368'b10010001000000010111011000010011010110010010111011010001101101100100000000010001011010001001101000001000011001010101100011001101111100010010101100010010111001011110110100101001001100111100011101011001010001010001111000110110111111010001100000001100010001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000101010000;
neuron_parameter[22] <= 368'b00000010000000000101110110001011100110001010101010001111110110101000111100000010010011111001011111001101101000101011100001001011001001100010001011010010001000000000001111010100001101001000011001001101001101000110100100101110101000001011011011001010110011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000101100000;
neuron_parameter[23] <= 368'b10101000110111101010111110101001101010010010101011101010001010110010001000101010100010101010101010101000101011101010001010101111101010101010001010100000100010101010001010001000100000101010101110001010101010100000100011100110101001001010100011001011001010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000101110000;
neuron_parameter[24] <= 368'b00010010000001000010101101101010100100000110001001100111100110101010111010010110010001100100010000110001000110100010010010100010011010011100110111101101100010000011010010100001001100010111110010111010101010110001011100010100010111101000000110000010000101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000110000000;
neuron_parameter[25] <= 368'b10100001110100011001001010011000010001000010000010001000010100011011011101101100100010110000111001001000110000000010000101000110010111110111010100011001110101110010111001100011100011101010110101001000000011001010000000101011000101000010011001010000000100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000110010000;
neuron_parameter[26] <= 368'b00101010100010000010000000011110110110100100101011001010101100100100110111011011010001110110001110010111011110001001011010111010011001101110000001001001000010101011101101110000110110011101101100001010111000110001010000110110011111000000110010111100001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000110100000;
neuron_parameter[27] <= 368'b00010100001101000010111111100110111100010000101100100111000010011010101110111110010001110100010111010011000101100011010010010001000001100000011000000001100001010101111000001110001101000000001100100100101111100110101110001100000000110000001111110001011101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000110110000;
neuron_parameter[28] <= 368'b10101011101010101010010010000011011000010010000000001000001110101101000011101010100000101110000010111110000110101101101101111111101110101110100100001010011000110100101010101111101010101011100100000001100000101111110001101001101000001110001011001010001011110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000111000000;
neuron_parameter[29] <= 368'b00110000000100000000101011100101111111010000100001000011100010110001101100001110011001100000110111111010001000100110000010110000100001101011011001000001001001100000101001000010110010001110001100100001001101001110100100100011010000010010111001111001111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000111010000;
neuron_parameter[30] <= 368'b00100010101011001000001000001110100001001101011001001010101001100011101111101010100000010011101110001111111011000011001000000010100000001001001001000101100011110110000000000110001010001011001010100101000000100101001100001100001000111010101010001001101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000111100000;
neuron_parameter[31] <= 368'b00010110001100011110111001100101110100001100110100100111101001000100000010111011000000001010000011010011001000001101101010101000011010001001101110110110011000001110000110001000000100101100000010101010111010101101111010110011100011100000000110001010100001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000000111110000;
neuron_parameter[32] <= 368'b00100011000010110111011000011001000011001000100011001110011101000100110101110011110001111011000000001101111000001001010010001110100000101000001001000100001011110000000001011000001111000000000000000001001000101100001000000010100000101101011110110101100100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001000000000;
neuron_parameter[33] <= 368'b10101001110111011100000000111001001001100011001010011000010100010111101001100110100100001100000000110001101000110110001100110111100010000000001010010100010000110101001000000111101101100010000001100100000000000110001001000111001000101110011110110011100110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001000010000;
neuron_parameter[34] <= 368'b00010000001100100111111111100001101100011010101000000101100010111000111010000110101100100011110111010000001001111100010011100001011010011100110100000100000011101011010001100001001000011111011001010110110110111101010010010100010111010001100000001001100000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001000100000;
neuron_parameter[35] <= 368'b10101001110010010000000000010000001001101111000001011000010001101111001100101000100110110110111001001000010000101010001101000101110111111101000110101010110101100100111001000001100110101100110111011010110110001010100010111001010011000110001000000010011110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001000110000;
neuron_parameter[36] <= 368'b01101010110010001000010001000000100100100000100100101010111100000111011111011001100000000101001110111110100010111001011010110110000101001111000010001010110111001011101001110000100110101000111011001010000010010011110010110010001111000010010010001110001000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001001000000;
neuron_parameter[37] <= 368'b01011000001001100000101101000110111100010001000000100101001010011010111000111100011011011000100000000001000111110010000000000011101110000001011000100100101010010101010010101101000111000001100110100110001100100010001110111100010111000001000110000010111101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001001010000;
neuron_parameter[38] <= 368'b00101111111011100000010100011011100001100101111110011010101101100101100111010001111000010101001110101110011110101101111011101111101101100110000100111011000110100100100011010111110000101001111111000001000001001111000001111010100010011110011000100011011000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001001100000;
neuron_parameter[39] <= 368'b01010010001100010010100010001000011101010000100000000100000000011001101000101100001111100000110000000000101001000010000101010001100100110001110101000101100010000011000000100010010010011011001000000101000100010000100101000001001000111110011001000101011010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001001110000;
neuron_parameter[40] <= 368'b10101111111010101110010010111001100000101011110110101000011100100101111101101010100010111010111000001001111111001001001111000010101001100000111000000111101010111011111110010010101000001111001001001001001011001110101010101010101010010000101000100000101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001010000000;
neuron_parameter[41] <= 368'b00111000101010000111101101001110110000011001011001100011101011000100000000110000001010000000101000000000110011010011100001001101110111001001100110011010011101001111101010011000001110101100011011011001000001010101110000011100101001001110110010001010001001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001010010000;
neuron_parameter[42] <= 368'b10000011000010110111110010011001000010100110001111111110011100100100110001010011110001011000000100101101111100101001100010001011000011100011001010010100001000011000001101011000001101000000000101100101000001100100001000001101101000101101101011010000101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001010100000;
neuron_parameter[43] <= 368'b10101001111110001001001010001001001001110011001000011000010100011011001000101110100110011001111000110100100010110110000100011111000000100011000000010110001001000101100110011011110001100110001000100001000000001110100011001000101000101100101001110000101111100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001010110000;
neuron_parameter[44] <= 368'b00011100001001100100100101000110111000010000010000100101000000001010001010001011011100000000000011111010000001101011100011111000001010011110100011001011000010100000000001111000001110010110111010000000111110111001111010110100010111111000000100101010000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001011000000;
neuron_parameter[45] <= 368'b11101101110110011000000000011000010001000010100001000000111001001111110100101000100101110100111001001001110001100000001101000100010111101111000000101011110101110011110001100101100011101000110110010000110111011011010011110001010010000010100000000110011110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001011010000;
neuron_parameter[46] <= 368'b00101010110011000000001100111110100001000110001001011010101110100111100111011011010000010110001110000001011100000010010000011110001011111111010001101001100001100001010001110000100110000010101010001010111010110011010010100010010111110001100000101110100000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001011100000;
neuron_parameter[47] <= 368'b00001110001101100111110001100110010110000110001100110111001010001010110010100011100001001000000111111011000111100001111000110100110001000000101010000000001000000100001110011101001100100000001100100000000000001000001111001010100000101110011100100001101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001011110000;
neuron_parameter[48] <= 368'b00101011111010101000110110011011001011010001010000001000000100000101011011101011100010100110011010110110111110111101101011110111101100101110100100101010001010010100101110101111001000101011100000010010000000001010010000101001011110000101011101111011001010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001100000000;
neuron_parameter[49] <= 368'b11010000000101001010110011100000011001010000000001000000010010101001101000000110000100100110111111110110101001011100011000010000110101100101100111010100001100101110100000011010001000011101110000000001000000100010101101000001000000111110111010100000101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001100010000;
neuron_parameter[50] <= 368'b10100110110011001000000000011000000011100101010101001000010100000111101101101000100010011000110000001100110011000011001101000110010100010011110100001110001101011110000110000011111000111111000001101010000000101110000000101110101000010110011011000111100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001100100000;
neuron_parameter[51] <= 368'b01010010001100000100101101000111110100000000000100100111101011010100000010101010010000000010000110010110000101110101100001101000111001010111100111110110010101001011000110111000001100111101010010110101111010111101111110010101110111100001100010001000100011110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001100110000;
neuron_parameter[52] <= 368'b00110010000100000101100000101001100110101100101011101110110110111010001111100110010011111101110001001001000100100011100011101011001011100000000011000010001000001000001101010001001101000000100010001101001001000100000000001000101000101101001011110010100111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001101000000;
neuron_parameter[53] <= 368'b10100000100010101011001010010000001010110011010000010000010110101011001000101100100010110000111001100000100010110000100100001101111100010010011110010010001100001110011110011101001000110000000010101101101111001000001010011100100010011000011001010000111001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001101010000;
neuron_parameter[54] <= 368'b00011100011000000100101100000010001110001010111001000111000011001011011110011110100100111101010001100000001100000000010010100000011110011101111011101111100011000101000001110001101110010101110010010010001000110001011011110000100101011110100100101010100001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001101100000;
neuron_parameter[55] <= 368'b11101111100110010000000000010010011001000011000100001000000000101101111101001100100000111100110101000000011110001010011101000100010111101111000001101001110101100001110001010110110011100010011000001001110111011011110011111001010010000100110000101110011110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001101110000;
neuron_parameter[56] <= 368'b00100010100110010010010100111000100110100101000011011010111110100111100111011001100001010100000110010111011111001101011010011110011100111110000001001000000000101011110100110000110110001110101001001010101000010010010000111011001111000001010010011000001110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001110000000;
neuron_parameter[57] <= 368'b10011000001000100011001101000110011000001101000000100111101010001010111010101111000101011101110011111110100011100001001000110000110001000100001010010010001100001100001110011101001101100000000110100011100000000010001101011011110010011010001110100001100100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001110010000;
neuron_parameter[58] <= 368'b10001111101010111000010010011001000001100000111110101010000101101111100000010011110000000110000110110010000011111101111010111001001000110010100100010011011000000100000111100011101000100110100000100100111000000010001000100010010000001000011000111100110110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001110100000;
neuron_parameter[59] <= 368'b10110001010110000000110010100001001011111001110000001101000011011001000001100100001110101000101000100100101001010010010110000010111000011000100101100101001110111100100000001010001001110111000001100000000000110000101101000010001000111110111110101011101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001110110000;
neuron_parameter[60] <= 368'b00100111111011101000000000001011001000100100011101111000101101100111111101101010100011110010111100000110010011001011001101000010101000101001111010000100101011110110110000000010001010001010101001111101101011110110101010001010010010110011101110001100111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001111000000;
neuron_parameter[61] <= 368'b00011000001100101110101101010111110110011101100000000111101011000000000010111001001010001010101010001110011000001011100001001100001101000111100010110010110111000011100111101110011010101101111111010111011000110001110001010101011111101111011111001000111001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001111010000;
neuron_parameter[62] <= 368'b10000110100010101010000010011010000000100001010110011010111111000000000011010001011001011000000001101101110111000011110000010011101001100000000100010010001000011100001110011101001101010000000101001101000011000110000110010100100010011101001001000100011111010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001111100000;
neuron_parameter[63] <= 368'b10101001111110001101101010010001001001000011000010001000010000010011001000101101100010001001001001110000100000110100100000111101100100100000011000010000000000000111001110001111100001100010000110100100010100100000001101001000100000101110011011110001101110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000001111110000;
neuron_parameter[64] <= 368'b00011010011110100100101110100000011011001000101010010100000011101010111110011010010001110001100011100001001001100010001010110000101000101010111010000010100010101011011110101010001010011000001010111101100000011101111101000111101110000100000101001100010110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010000000000;
neuron_parameter[65] <= 368'b10100010100000010000000000011000010010101110011110111010111100001011000000001100101110001001110000101000110011010010000100000101110111101101100111101011110101101100101000110101100110101100010111001010000011001010100010100001101000000110011000110111010110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010000010000;
neuron_parameter[66] <= 368'b10111010011010111000010000011000100001001000110000011010101100000111111101001000100000110111001000101000110010101001101010000010011101001010000100001010110111001010101011100001100010101000011010001000100010001010100010110010110111000001100000001100000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010000100000;
neuron_parameter[67] <= 368'b01010000011100001100101010000100100001010000110000000100100010011111111001101000001110100010110000000000110111100010000101000011100010111011011101100001100011011011010011100010100011011010010010011010100010110000010010001001000011100011101010011010101110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010000110000;
neuron_parameter[68] <= 368'b00101110101010101000011100000000100001101101011010001001100100000000000010011001011100001111000010100010011010111101100011101111000010101000101001101001001000110000000111000110011010001010010110110000001101001010100111110000100010001101101100101111011010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010001000000;
neuron_parameter[69] <= 368'b00010010000101000100101101100100111010010000000011101111110010111001101100011110011100100101110111111010001001001100011010110000000001100101100100000000010001100010100001100010110010001111101100001000100111000110100110001001101000010010101011110100111011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010001010000;
neuron_parameter[70] <= 368'b10101101111010101010000000011000000010101101110100101000101001100101111101101010100010010010001100001111111011001011001101000010111110110101011000000011101110110111010010000010110010011111010000100001000001100010001100001011011100111011100010000001000011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010001100000;
neuron_parameter[71] <= 368'b00000111011100111110110001100101110100000100111100100111001001000000000011111011000000001010100010010011001000101111001010101000101010001000101110100100011000001100001110001100001000101100000000101010111011101111001010100111110111101001000111001100100101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010001110000;
neuron_parameter[72] <= 368'b10000111101010101011001010001010000000100001110110011111111110100000000011010001011001010101000001111111110111100001110010111011101010100010000000010010001000111000001110011101001101010000000100000101000001000110001101000001101000111101001001100000110111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010010000000;
neuron_parameter[73] <= 368'b10101101110010111001000010001000001001101101010101101000000000011011001000111100001110101001101001101000100010000010000100000101111101010010111100011010100010001011000111011001010101110110100011100110001001000100001101000110101000101101010010100011100101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010010010000;
neuron_parameter[74] <= 368'b10011000000110000110101111100001011100011000000000100111100001001001110010010111011100001101110111110000000111010000010010100000111010001110110100000011100010101011000010101001001010011101111011011110110010101101111010010110010111011000000100001000100001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010010100000;
neuron_parameter[75] <= 368'b10000100111100101001101100001100011001111101000001000100110010010110000110100000111100110011101111101100111000011100010010101000101110111010000000111101010011111111011100101010101001110010000110111110111100110000001110000000001011100001101011011010111110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010010110000;
neuron_parameter[76] <= 368'b00101010100010000010101001101110110010101110001001001010111000100010100111011011010000010010101010000010011111000000000001101010000011101111110011101000000000101011101000110000100110011101101011011010010000110001011001110110011101100110010010011110001000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010011000000;
neuron_parameter[77] <= 368'b00011000001101100001100011100110111100011000100100100101000010010010100110011111010000110100010111110011001101100011000010110000100011100011011000000001100011010001011000000110111111000000001100100000111100010100001110001100000000110000001110111001111101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010011010000;
neuron_parameter[78] <= 368'b00100100100010101010111010101010101010111010101010101000101010110000101010001111011100101010101010001010101010101010100010111010101010101010101010101010101010111110001010101110110010101010101001101111001000010110001010111000111011101000101000101011101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010011100000;
neuron_parameter[79] <= 368'b10101010100100100011110010101010101110101000100011001000101111001011101111101110110011111110111010101010101110001010011010101110001010001011111000100001101010010001100000100010111010111001000010101010101010001010100010101010101010101010101010101010101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010011110000;
neuron_parameter[80] <= 368'b00101010111000100010101010101010111010111010101010001100101110101010110010101010101110101010101010011000101010101010100010000010101010101000100010100010101011101010101011001010001110101010101110101000001000101110111010001110111010111110101000001010001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010100000000;
neuron_parameter[81] <= 368'b00100010101000110011011010000111000110000011000000011011001010000000000000010101011110001001101000001100111110010011100001001101010000000001100110010010111101011111101000001001000100111000000101111000001011100101111000110110111111010000100000001000110001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010100010000;
neuron_parameter[82] <= 368'b10100010100010000110010010101001100110101000101111111010111100100010011001010110100001111101001000100001000110100000100010101011100001000000000001000000001000011000001010001100001111000000010110100101001000100000000100000001100000101111001011110011100011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010100100000;
neuron_parameter[83] <= 368'b11100001110111011101000010110000000001100011001100001000010100010111001011000001100000001101011000110000001100110100100000111101100100000010000100010010011000011110001110001111000001101000000100100101100001100000101110001000100000101001010011110101100111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010100110000;
neuron_parameter[84] <= 368'b00010001000010000110111011100011010000011010101000000111101010111011011010001010111101100000110011110000000001001010011110100000101010011010101011100111000011101001000001110010001110010111011000011010110000111101111000110110110111011001000100001000100001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010101000000;
neuron_parameter[85] <= 368'b01101001110010011001000000011000000001101101110010011000110101010101001101100010100100100110011111100100110000101101101100100101111101000101001110011010110100001010111111001001000001111000000011000010000000001010100010101110010110001110001100000000001000110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010101010000;
neuron_parameter[86] <= 368'b01101010100010111000000000011000100000100001010011011010001100000010000001011001000000011001001000101000110010000101011010011110000101101111000110101010010101100010101000110000100010101000111101001000000000010011010001010010011101000110010010011100000000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010101100000;
neuron_parameter[87] <= 368'b10001101001101101110110111000010011110100100001110100111001000001100111010101011000101001000010011110011000101101011111010110000100011000000001010010010001000101100001110011100001100100100001100100100100100000010001111001000100000101010011110100011001110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010101110000;
neuron_parameter[88] <= 368'b00101001111010101000010000000011001001110001010000001001000010000010011100010010111001100111101110100110000100110000100001101001001110110111100001101001100110000000100111110011010000001011111000000001000000000001000011010000000001011110111100000000000000110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010110000000;
neuron_parameter[89] <= 368'b01010010010101100100100011101100111101010000100010100101010010111001101100111110011100100100101111111110101011010010000110110000000000101101110101000111001011101100100000100010111010011111000000100000000101100110101110100010101000111110101010100111101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010110010000;
neuron_parameter[90] <= 368'b10100101110011111100011000011010000010100100011101111000111100100111111101101010100011110011011100000111111011001011001100000010110010011001011001000001100011110111010000000010000010011011001001010101000000100110011111011010001000010011001011001000001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010110100000;
neuron_parameter[91] <= 368'b01011010001100101110111101100110001100001100000100100111101001000100000010101011000000001010001110000011001000000111101000101000111000001000101110010110011100001110001110001000000000111001010010110101111011100101111010010101111111010001000110001100010001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010110110000;
neuron_parameter[92] <= 368'b00100110100010000100100010101011101101101011001100111111010110111010111111000110110001111101010000100001000110100010100001100111000011100000001011000000001000101000001001000000001101000000111001100111001000000100000000001100101000101001001010101101110011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010111000000;
neuron_parameter[93] <= 368'b00101011010111011000000000010000000000000100001011001000000000000000000000000011100000001101000010110111001000110100100000011101010100010110010100011010011100010111010110101001010001101000000100001101100011000100100010011000000100010001100011000100111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010111010000;
neuron_parameter[94] <= 368'b10010000000000000111101001100011011100000010101001100101101000111000111110011010111101101001110101110001001101000001011010100000001010011110110111100101100011100001000001110001001110010101111010010010111010111001011000010100010111011000000100101000100001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010111100000;
neuron_parameter[95] <= 368'b00000110000000000001100100111000100000000100001011100010110110101010100111000000101001110000101111111000111001111100010111001011111011111001000000100011110100101010011100001011100000100010000100010100111110110000001110000001000010101001101010010000110010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000010111110000;
neuron_parameter[96] <= 368'b10100010100011000000000100111000100010100000001101111010001100111010101011111111010010101000101010000011001110001110001100001010000011101010111011001101000001101100110000101000100110000111101011011000001000010001111001000111011101100110010110011110000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011000000000;
neuron_parameter[97] <= 368'b01010111001100001110110101100110110010011100010100100101000000111101110011111100011011011000000000000001100010000010000110000011100100010100001000011000101101010110111010001001001001100000000100000000110110101010001101000011000000001110011100100000101100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011000010000;
neuron_parameter[98] <= 368'b11101111111010110000110100011001000100100100111110101000100001100100000010011011111000001110000110110010011100111101111010111101000000101110101111101101011000100100000110111011111000100011110000100101001000111111011001000111010000011011010100101110101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011000100000;
neuron_parameter[99] <= 368'b10011010000110101101111111101010011000101000001010100000100011001000111010101000101110111010111010101000001010101010101010101011101000101010101010001010000011011000001000111100000010101010100000111110011010101100000110000010001111101011101111100010011010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011000110000;
neuron_parameter[100] <= 368'b10101111110010101000010000111011000000100001010111111000100101100111101101101011100011110011011100001111111011001011001001011010110010101001011001010101010011110110110000010010101000001011001001101101000001100101010111010001001011010011101010001001001011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011001000000;
neuron_parameter[101] <= 368'b00000010100000000111011100000011000110000011000001001011001110000000000000010100001010001000101000001000110111010010100001001101100000010010100100000010100001100010001000101010001011101000111111010101010000110000011001000100011001000101110010001010100010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011001010000;
neuron_parameter[102] <= 368'b00100010100000000111110010101111100111100010001111111110011110110010111011000110100001111101010001101010001110101010100000100011000011100000001011000000001000101000001001001100001111000000001001000101001001000100000000001101101100101101001010110111100111000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011001100000;
neuron_parameter[103] <= 368'b11001000111111001101101010010010001011000010000000001000010000010010000110101111010000001101101001110110101000110100100000111000100011000000001010010000000000001101001010011101001001100000001101100010001100100010101111100010000000011110001110110010100010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011001110000;
neuron_parameter[104] <= 368'b00011000001000101101011001000111010000010011001000000101000011101000101010000110101110100110110110111010001101110000011111010000001010111000110100110101100011001011010111100001000000011011011001011101110011111111110010111100010111010001000001000100110001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011010000000;
neuron_parameter[105] <= 368'b10101010110110000000001000001000001001100100010000011000010000000010001000101010000110001000001001000000100000110010100100000101010111101111100011101001110101100000100000110011110010100100110110010010000110001010000000100001010010100010000010101011010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011010010000;
neuron_parameter[106] <= 368'b10100100100010010010001000011110100000100000011000001010001000100111110101011010000000110000101010001001011110001010001001001110000111011111000011001011000011100011101001110000100010001010111001001010011000010001010000110010011111000010010110011110000100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011010100000;
neuron_parameter[107] <= 368'b01011000001100101100100001010110111000010000100100100101000000011001111001101000001010101000100000000001100011100010000111000011100010101000011001100000000011110011010000000110110011000010000110010000001100110001011000111001000010000000001110101000001100010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011010110000;
neuron_parameter[108] <= 368'b01101110001010110010010101011000110000100100111110100000100001000100000010010011011000000100000110100010000100101101110010101000001000010110101111100111011000101100000111010001001000111001100001100010001010101010001010000010000000011001001101110001100000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011011000000;
neuron_parameter[109] <= 368'b00000000000101000011001001010001000101010000001001001100010000101011011100000110100100100110110111110010000010100000000000110100011101010111101110010010011100001110000110010001001000110101000000100001000011000010101111001000100000011010011100010000111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011011010000;
neuron_parameter[110] <= 368'b01100110111011101000000000001010101001101100011101101010100001100101111111101010100011010000110110001111011111001011011101000010101000111001000000010000100011110111000010000010000010011010001000001001000011101110101011010000000010010001101000001000111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011011100000;
neuron_parameter[111] <= 368'b10100011001000110011111110001011000111000011010001010001001110100100000001010101011010001001101010001000111100010101100001001101011000000001000100010010111101010110100110101011000001111001000011101010111001010101011000110110111111000001000000001110010101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011011110000;
neuron_parameter[112] <= 368'b10000111000010010011010010011001000010100100101111111010011100100000100011000011111001101001000000111111111100001101111010001010000000100011001100010010001000011100011100001100001101001000000100001101100011100100001001101010100000101001001001110000110010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011100000000;
neuron_parameter[113] <= 368'b11100001111011101000001000110000010000110011001001000000010100111011001000101100100110001000111001100000000010110010000100001101100001000010101010010010000000001000000110011101100000100100001100100100001101101100001000001110100000101001011111110001111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011100010000;
neuron_parameter[114] <= 368'b00010100001100000111100101111100011100010000010110110100000001111010111010011010110100101001000110111010000011100000001010101000101100011110101000011110100010001011001110111010111110111100100010011001000010011001111011010000101010111100001100001000001000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011100100000;
neuron_parameter[115] <= 368'b11100111110011001011001010000010111000011001010011100000110100011010000000000000001100000001011011101000010000010010100000100101010111111111000110101011110101100110111000110001110110101000110100000010100110011010010010101001000000000010101100111011010010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011100110000;
neuron_parameter[116] <= 368'b10100010100011000010101001101110111000000110001001111010001110100010001011011011010000001000001000100011001110000110000101011010000001001111110011001000001000101100100000111100100110001111101111110000001000110001110000010110011101100010010010011110001000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011101000000;
neuron_parameter[117] <= 368'b00011000001000000111110011000010111000010000100110100100001000011001111011111101011011011000000000001001000111000011000110000011100000000000011001000100000011010101011000001111001011000011000110110010111100101010011110001001010010100000101111111000001101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011101010000;
neuron_parameter[118] <= 368'b10101101100010101010000000000010000000110011001110101010111110100000000010001011111011001110001010111110101100011101111011111100000110101010000000101000011000100001110001100100110010001010111100000000000100010111100111001000001010010111101001100111011011110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011101100000;
neuron_parameter[119] <= 368'b00010100000100001010100101001010010000010000001001100110010011101001011100100110000101100110110111110010001001000010010001010000011100010111100111011101011110001110100110110010111000110111100001010001000000101000101001000110000000111110011100010001101010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011101110000;
neuron_parameter[120] <= 368'b10100101100011011000110010001010001010100010110110111000010100000111111101111000100010110010011000000000111011001010001101000010001010111001000000110001110011100111100011010010100000001000011010001011101000101010001000101010111100010011100011101100110001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011110000000;
neuron_parameter[121] <= 368'b10010010000100010110111100100100110000010100000101101111111010100000000010010001000010000000000011010000001101010011100001001000101000010101110110110100111100011111110110101000000100111101010010010110111010110101011110000100110111100001100010001100110001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011110010000;
neuron_parameter[122] <= 368'b00000011000010010110010000111001100110001100100111111010111100000100000011000011110000001010000011111111111100001101111010001000100000000000000100010000001000011000001110000101001001001000000100100101100001001110001100100001100000101011101011110110011011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011110100000;
neuron_parameter[123] <= 368'b10100100110010011010001000101000100000100011000101111000010100010001001100101100001110000001100001101000000000110010000100001100111100010010111100010010010010000110001111010111111000110110001010101111001011001100001101001010100000101101001110100001100110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011110110000;
neuron_parameter[124] <= 368'b00010000000001000110111101100010001110000000101001000111001010011000111010001110011000101001110001110010001100000000110010110010001010111000100011000101000011101001000000110001001110010111111011010000100000111001011001110111100100011110100100000011100000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011111000000;
neuron_parameter[125] <= 368'b10101001111110011000001000001000010001001010000000001000010100111111110100101000100010111001111001001000111000100000001101000110010111111111000100101011110101100001111001100111110011101000110100001000110101011010010000010000010111000000111000010100010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011111010000;
neuron_parameter[126] <= 368'b10100010100011000000100101111000100100000010001101011010001110110010001011011111010000001000000010001110000110010010001001001010000101001111110011001000001001101010100000110000100110101100101011011010001000010001110000110010011111000010010010011110001000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011111100000;
neuron_parameter[127] <= 368'b00011100001100001010010011100110111110111101000110100111101000100000100010010001001010000000000011101010000110000011110010001010100000000000011000000001001001011110111000001101001001100000000100100100110100101110001010001100000100110010100000100001111110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000011111110000;
neuron_parameter[128] <= 368'b01101110111011110000010100001001100001001100111110001010101000000100000010011011111000001110001010100010010000101100111011101111000000101110000001101101001000000000100001110011111010000011110110010100000110011010110001101000111000011110101110101011000010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100000000000;
neuron_parameter[129] <= 368'b00111000001111001010101011100110111100010000001010111101101010101001101010001111001101100100100111111110000001100110000100110000000001100010110000000000101001100000101001100010110000000110101100101111011011101110100010101110010110000001101001010101111011110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100000010000;
neuron_parameter[130] <= 368'b00101111100010101010010000011001000000100101011100101010101001100111111111101010100011110010110110000111011011001011001101000010100010001001000001000101100011100111010000000010110010011011001001000100000010110100111011010011101110111010101000000010001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100000100000;
neuron_parameter[131] <= 368'b00010011001100000110110100100111100110000100001001101111011010100100000010100000001010001010001110001101011100000111000001001000111011010001100110110010111101001111101110001100000110111100010110010111011010110001111100010101011111110001100010001000010001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100000110000;
neuron_parameter[132] <= 368'b01101010100010110010001000011000000001001000110010001000001101000100000011110011011010001010000000101101111000001011011010000000100000000000000000000000000001001000001000001100001010101000000100100000000000100000001101000010100000101101011110110011001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100001000000;
neuron_parameter[133] <= 368'b11101101010111111100000110100000001001000010000111001000000000011011101100111100010010011001110001101000000010001010000100000010111100010010111100011010110010010011000111111011000111101010100110101110001010000100001100000110100000101101010110100001100101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100001010000;
neuron_parameter[134] <= 368'b00010100001000000101111001100100010100010000000000100101000010101000111010000100001111101010010100110001001001100000010111110000001010111000110100100101100010100000010111100001000100011011110010111010111010111111011000111100010111010001000101001000100001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100001100000;
neuron_parameter[135] <= 368'b01100001110000000001001000010000000001100101010001001000010010011011000000101000100010101000111001101000110000010000000101000101010111101111000100101011110101100000111000000001110110100100110110000010110110001010000010101000000000000010001100010001010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100001110000;
neuron_parameter[136] <= 368'b10100010100011000010000100101010100001100110001101011010111110110010000011011001010000011000101010001010100110010000001000111110000110001111110010001001011011001011101000110000100110111100101011011010011000110001110000010110010111100010000110011110000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100010000000;
neuron_parameter[137] <= 368'b00011100001101000010100111100110111100011001001100100101000010000010110010111100010011010000000000000001000111100011000010000011100000000000011000000100000001010111111000001110000111000001100100100000001110101010001110001011110010100010000110101011101100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100010010000;
neuron_parameter[138] <= 368'b00101111111010100001010100011001100011001000110110001000000000000100010000011001011010000111001110100010000100111100111011101101001110111111001101101101010011110000100001000011110100100011110010001010000100001011000100101010101000101010001100110011000100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100010100000;
neuron_parameter[139] <= 368'b01011100001101001101100011000110011000011001000010100101000010001000000001001010011100001010101010111110000001001110000110110000000100110000110100011000001010100010100010100010110010111111100000100010000111100010101110001001101010110010101011010101111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100010110000;
neuron_parameter[140] <= 368'b00101101110010101000010000011011001001101110011100001010100000100101111111101001100001110011011110001111111111001011001011100010101011100001010001010101101011110010110001010010010000011010001001001101000001100100001100001000010010110011100101100100110011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100011000000;
neuron_parameter[141] <= 368'b00010001100100010111111110000011010110000010000001000101010010000100010000110101001010000010101001001100100000010010100001001100100010001000001001010000011001010101001000001100000111100000011111011100011000110001010000100101111111000101010010001010110000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100011010000;
neuron_parameter[142] <= 368'b10000010001000010111100010001001000111001010001010011110001010100100000101100010100000111011010111101101111000101011101000100110001011100011001001010010001000001001001101011100101101000000001101001101000000000110000000101110101000101110011010000001100001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100011100000;
neuron_parameter[143] <= 368'b11001000110010011001101000111000101001110111010000000000010000011011001100111100101110000001111001101000110000100000000100001101111101000010111110010010010000001111001110011001101101110000001000100100001010000000001100001010101000101101010010100011100101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100011110000;
neuron_parameter[144] <= 368'b00010010000001000111111101100110000110100110001001010100100100101011011010011110011101001000010100100000000010100011010010100000001010011110111111100111000010000001010010110000001100010101111011011010001000011001011000010111010111001001000100001010000101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100100000000;
neuron_parameter[145] <= 368'b11100101110110011000001000011000010011001101110011001000110001010101000100100000100100000100111011011100100000000001101001000111010101100101000100011010110101110010111011101001100111101000110111010010110010010000000010011001001010000110011000000010001110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100100010000;
neuron_parameter[146] <= 368'b01101110100010110010001000111010100010100101010001111010101101100010001001011001000000011101001000101000011110001100111010011110010101001110000010001010010000101010101000111000110110101000111101000000000000010000010001010111010101000110010110011100000010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100100100000;
neuron_parameter[147] <= 368'b00010110000101000010100101100110110110010100001101100111101010101111111111111100011011011000010000000001000110000011000111001011100000000000001000010000000001011101011010001101001101000001000110100001111101101110001101001101000000010001001000100100111101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100100110000;
neuron_parameter[148] <= 368'b11101110111011101000000000000011001010101000110110101000101101101101111010001011110000101110000010010011000110101101101011110101100010111110000101011001001000010100000111111010001010101011110101000001000000000010110101001000001000001100011100101010000010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100101000000;
neuron_parameter[149] <= 368'b01010000001101000000101100100100011010010010100000000100010010011001101100101110001111100010110001100000000001000010000101010001101000111000110101001101101110001000100001100010110010010111010000100001000110101110100111000110100000111110011001000001111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100101010000;
neuron_parameter[150] <= 368'b10100101100010101010010010101011001010100010010011111000110100100110111001111000101011110010001000000110111011001010000000010010011010110001110000010000001010100010010111010010100010001010101011001100101011101110101010001010111010110011100011011000111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100101100000;
neuron_parameter[151] <= 368'b00010000001100010111011110000111100100001110110001000111111010000000000010111100101010001010101000001000111000010011100001001100001101001011101110101000100111010111100010101010000010101000111111110101011000100001111000010100001100101111111011001010011001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100101110000;
neuron_parameter[152] <= 368'b10000011100010110011000000011000000011000000110011011110011101010000100011000000011011111000000001101101111010101011101010000010100001100001011010010010101000011000001100011100001101000000000101000101000001000110000001000010101000111101011011000000100011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100110000000;
neuron_parameter[153] <= 368'b11001000111100111100101010011000011001111010000000100000010000010000000100101100101110000001111001101000100000110000100000101101101001000010001010010010000000001110001111011101101100110100001110000010000000100010001111001010100000101100011110100001101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100110010000;
neuron_parameter[154] <= 368'b10011000000100000111101100110011010100010000100001110100101001101011111110010010010101101101010011100000001111100000001010100000101110011110110100111110100010101011011111111000000110011001011010011001110010110001111011010000101010111100001100000000000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100110100000;
neuron_parameter[155] <= 368'b11101001110000000000101010000000011001011111110001000000010010000010000000100000100100000011001101101000100000110010100100101100010111101111000001101001110101100000101001010011110111100110110110100010101110000010101110101000000010000010101000111001010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100110110000;
neuron_parameter[156] <= 368'b00101010100010111010000000011100100010100001010001011010001100100010001001011001000000011101001000001001110110000011000001001110010101101111000010011000000100101010101000111000110110101000111011101000000000000000010001010011011101000110010010010000000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100111000000;
neuron_parameter[157] <= 368'b01011110001101001011110011011010011110101010101100100101000000010110101010111001000010011000000100011001000101100101001110000110000001101000011000101001001010010101111010001111101001000000000110100110111010001010001000101001010010100010001110111000101100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100111010000;
neuron_parameter[158] <= 368'b00101110111010100000010100011001100001000101011110001010000001000111010100010000101000010111001110100010110010101000111011101111000100111011000000110001110110100010000101010010110010001011111000011001000000010001111000011001100000011010011000000100000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100111100000;
neuron_parameter[159] <= 368'b10010000000100100001110010100000101111001000100011000111100011011011101110000110011000111010100110110110101000101110011000100010101000101000101011001001001010010100100000001010111010101111000000100000001100110010101100000000101000111110101110101010101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000100111110000;
neuron_parameter[160] <= 368'b10101111111011101000000000011100001011100101011111001000101100000111111101101000100011110010111000000110110011001011001000000010101010101001101000110001101011110111100001010010100010001010001011001101000011101111111011001010001000010010101000000001101001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101000000000;
neuron_parameter[161] <= 368'b00010001001100110110111100000011110000011010101000000111101010000100000010111101000010001110001110001100011100001011100001001100101000000011101110011010111101000111101010111100001010101000011001010111001000110001111010010101011011101001100010001000110011010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101000010000;
neuron_parameter[162] <= 368'b00000010000000010111110010001011100010100010001011011110011110110010010001110110100001111111000001101101111110101010100000101111000001100001001010110000001010110000001101010000000101010000000010101111001001100110000000001011101000101101101010110010100110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101000100000;
neuron_parameter[163] <= 368'b10001000110010111001001010101000011001110010000110100000000000011011001100101100101110000001111001101000110000110010000100001101111001000010111110010010010000001110001111011101001100110110001000100100001001101100001001000010100000001001000010110001100000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101000110000;
neuron_parameter[164] <= 368'b10011000001101100101111101100011010101001000000000100111100001111011011110011010011110101100110011111010000001101010000011100000001010011000101011100001000010101011000001100000001110010111011010111110111010101001011010110110010111011000000100001010000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101001000000;
neuron_parameter[165] <= 368'b00000000100000001010101010110000000000100010001010101000010010100011000000000000001010010001111000101000110000010100110111101111110111111111000100111011111100111110111110001001000010101000010100000011111110010010010010001001000010011010101010000000001010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101001010000;
neuron_parameter[166] <= 368'b00100011110110000001010101111110100100000100101011101000101010100010100111011011010000110100111110010011011101001000010010111010011100001111000001001101000011000011100001110000110110000101101010101010111010111001010010100010010111110001100010011110000101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101001100000;
neuron_parameter[167] <= 368'b01011000001101000010000101100110111100011010001100100101001000101100110010111101011011011000100000000001000111000001010111000011110001000000011100001000001101011111111110001101001001100000000110100001000111101000001011101000100000101010001010000101111100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101001110000;
neuron_parameter[168] <= 368'b01101001111010100000000000001011100001000101011000001000000110000111010110111001110000011111001110100010011110101000101001101110001111101110000001101101100010110000100001010110110000001011111100000001000010001010000001000000100010011110111000110101011010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101010000000;
neuron_parameter[169] <= 368'b00010000000101000000111101100110011101010011000011000101000010011000001100011110001100100110110111111110000001010010010011110001000001100000100101101001001000100000100000100010110010011110000000000000000101000110101111101000100000010010101011111110101010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101010010000;
neuron_parameter[170] <= 368'b10100111101011101000000000011000000011100101010110011000110100100111111101101010100010010010111000001101111010001111001101000010111110011000101100010010011100010111110100000010011000111111000001101000000000100010000001001011101000101110010011001011100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101010100000;
neuron_parameter[171] <= 368'b00100101011100001110110001100101100000001000010100000111101011000100000011110001000000001000000010011011001000000101100010111000111010001001101010010110011000001110000110001100001000111000000010110001111010100001111010110010101011101000000010101000100000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101010110000;
neuron_parameter[172] <= 368'b00100011100010110111010000011001000100001001110111011010111111000100110001110001100011011000000000111101111000001101011110001110100000100001011000100101101001111100000000000100001101000010000110000101000010100000001101001010101000101101011011110001101100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101011000000;
neuron_parameter[173] <= 368'b10100010111010110000101010001011101010101010101011101010111110101010101010101010001110101010111010101010101010111011101010101110101011101010001100101000101010101010101110001110101011101010101010101010111110101000101100011001011011000010101011111011001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101011010000;
neuron_parameter[174] <= 368'b01011101001001100110010001100111011000011100000000100011100000001000011110000110011101001010100010101010000010100010000010100000001010111110100011101101000010100001000000111010101110000011111000010000111010111001011011010100111101111001100000101010000001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101011100000;
neuron_parameter[175] <= 368'b11100100110000001000100000011000011000001000110010100100110000010110000100101000001110100010101001001000110001001000111111101001111110111011011001101101110111110101010000101010101001110010000010111110001100110001001110000110000000100000101110010010000100010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101011110000;
neuron_parameter[176] <= 368'b01101110100011001010000001011110110000100001011011101010101011100011100111011001010000110110011110100011010111100000011000011110010110001110010010001000010010001011001001110000100110011100101010001010100010110001010010010010010111000010010010011110100000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101100000000;
neuron_parameter[177] <= 368'b00011000001101100000101100000110110011001010100000000101000010011001101001101100001011101010100000000000110010110010000101000011100010101001011001100001000011110101110010101010000011000000100110010010001101110111001100010001011010100010000111000100001101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101100010000;
neuron_parameter[178] <= 368'b00111110001010100010001101011111111000111101111110100000101000000010001010010111011001100110001110110010000111110000110010111001001100010100100110101111001010000000000111110011011000111111100001000100100000101000101010000010010100011100000100100000101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101100100000;
neuron_parameter[179] <= 368'b10010000000100001000110010101100111101111000100001100101000010011001001000001010001110100000101110111010001001011110001110110000101000101000100111000101001010110010100000101010011010011111010000101000000101101010101011001000100000011110101011110101111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101100110000;
neuron_parameter[180] <= 368'b00100111111011101011000001010101001001001100001100101000101001100111110111001001110001110001010110001111011111001011011011100010100011111001010000110101100011110011011001000110010000001010001100000101101011100100001010001101011010010011100011100100010011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101101000000;
neuron_parameter[181] <= 368'b00010010001000010111111110010111101110010011001100000111101011000000000010010111011010001001101010001011110101010101100011101100101000000000111110010100111101011110101010001101001000110000000111110100010001110101101000010100100001100100110000000000010001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101101010000;
neuron_parameter[182] <= 368'b10100000100010010111010010101011100110101011101011111010011100100010010011010110111000011101001001101001101110100010100010101111100000000000011000110100100010010000000000001100000011001000110100100111101000101010001000000010100010101010101110100001111010010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101101100000;
neuron_parameter[183] <= 368'b10111100101010111010101010101010101111101010101010101000001010111011001010101010011010101000101010101010101011011011101010101010101010101010101010101010101011101010001010101000001110101010000000000010111010101010101000101010101010101011101111011110111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101101110000;
neuron_parameter[184] <= 368'b00011000001100100100110111010111010100011000010000000101000000011011011010010011011101001000110011101010000011001011000000110000001010011110100011100101000010100001000000111000001110001111111010011110111010111001111010010110001111111001000100001010100001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101110000000;
neuron_parameter[185] <= 368'b10000100110011001000001010000010010000100011010001011000010100111011000000000000001100001001101011111010010000010010100100100101010111110111000100101011110101110110111000001011110010101010010100001010110010011010010010100001001001000010101000011010000010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101110010000;
neuron_parameter[186] <= 368'b00100010100001000011101100111110100111100100001001011010001110100111101101001011100001010111001110010101011111001000011000011110001011111111000001100001000000101001010001110000110110000110101011001011111011011011010010110010001111000001110000001000000100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101110100000;
neuron_parameter[187] <= 368'b01010000011101001100100001110100011100010000110100100101000000011001111011101000001011110010000000001001000100000011000101000011100010111001011001100001000011010111110011100010111011000010000100011110110100111000001000000001001010100000001110011100011101010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101110110000;
neuron_parameter[188] <= 368'b00101110011010100000000100011011100000011100110100101000101011100010011110010000111001110111001110110010010101111000110011111001001110010111100101101101101110000010000111110011010000011111110000000001100001110000111010100000100100011010001001001100101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101111000000;
neuron_parameter[189] <= 368'b11010000011100000010110111101000011101010000101000100000101011001001101000000100001111101000110010100010101011010010010110110000101100011001111101000101101010001110100000100010010000001111001000100101000001001001101111001000101000111110011000000101111010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101111010000;
neuron_parameter[190] <= 368'b10100111100011101000001010101001001000100010010111011000010100100111111101101000100011110010011000000110110011001011001101000010001011101001001000110001101001110010101001010010100000001010001011101111000001001111001001101010001100010011110110011000101011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101111100000;
neuron_parameter[191] <= 368'b00001111011100101110111001100101110100001100011000100111101011000000000010111100010100001010100010001111001000001111101010101100111000001000101110100100011100001100001010001100001000111100000001111110011011001101001010100100111111000001010111001100100001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000101111110000;
neuron_parameter[192] <= 368'b10100010000100000111110010001001001111101010101111101110010110111010111011000110110001111101000001111001001110101010100001101111000011100000000011100000001000010001001001010000010101000000001001001110000000000110100000001100101100001001001010100110110100100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000000000;
neuron_parameter[193] <= 368'b10101001111100001001001010011000001001100011001010011000010010011011001000001100100110001101111001110110110010110110100100001101110000110000011100011010011000010111010110001011110001110010001100100101011001101010100111001000101010111111101011010001101001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000010000;
neuron_parameter[194] <= 368'b00011100000101100110011101110111010100001110100000000111100011101001111010010110011100100001110111100000000001010010011110100001111010011000100011100110000011101010000001100001001110010101111001010000000010111001110001110100100101011100010100001011000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000100000;
neuron_parameter[195] <= 368'b00000010110100100000101000000000000001000010010000001000010010010011000000100000100010000000111001100000110000110000000000000101010111111111000100101011110101110010111000110001110111101000010110000010110110101010010110100001000000100010001000010011011110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110000110000;
neuron_parameter[196] <= 368'b01101110101010101010110000011000100110000100011101101010001001100111111111011011010000110100111010100001001111000010100000011110011110001110010011101001000010001011100001110000100110011100101010101010110000110000011000100111011111000110010000110000000100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001000000;
neuron_parameter[197] <= 368'b01011110001101000010010101100110110100111000001100110111001000101010010010111101110011001000000011011001000101000001100100000000110001000000001010010000001000011100011110001101001101100000001110110011111001001110001100100011110000110000000100100000110101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001010000;
neuron_parameter[198] <= 368'b00101110111010100000000100011000100001000001111110001000101101000110000000010001011000000111001110100010011110111100111011101010001000111110001101111101011010100100101011000010111000000011111011100010100001110010100000110010101000111010001001100100011010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001100000;
neuron_parameter[199] <= 368'b01010010000001001010101001100111011100010100000001000100011010111001101100100110000101100000110101110010101001010010010000010000001010110110100101000101001010101110000000111010011000010111010000000000000000110010001101000000000000011111111110101010001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110001110000;
neuron_parameter[200] <= 368'b10100001101010011000000010101011001000100010000110111000010100000111111001111000100010111010111000001000111010001010001101000010001000101001000000000001100011110011101001010010100000001000001010001001101000111011100000011000111000010011100110110000010011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010000000;
neuron_parameter[201] <= 368'b10010001001100010111010010010111000100010011110000010001001111000000000010010101111010001001101000001000101100000111100011001100100000000000100100010000111001111110101010001101000011101000010101010010001001110001110000011100111111010101000000001100111000000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010010000;
neuron_parameter[202] <= 368'b11000010100010100010001000001000100011001000110001001111001001100110100011110001110011011010000000101101111011100001110010001010100101000011001001000110101000111000001001011000100111000000010101100101000001101100000101000111101000111111011011100001000110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010100000;
neuron_parameter[203] <= 368'b10101000110101001101001010111001001001110010001001011000010110010010000000000100100010011001011000110100101010110100100000101101101000000000011000010100010000000100001110001111001001100000000110100110000111100100001101001110100100101001011011110001100101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110010110000;
neuron_parameter[204] <= 368'b00011010001000100110101000100111111010010010001000110111000010001011110110011010110001110001110111101001001110100010001010100010101000001000110000000010100010101011010001101000001110011010011011011001100000010001110000000000011010001100000100001110000000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011000000;
neuron_parameter[205] <= 368'b00000100110100001001101101101100111001010100100011100101110010110110000100100000001000100011101111101000111001000100111010101001101110111010001110101101010010111110010100101011101001110010000000111110111000010000001010000001000011100001101011011010110010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011010000;
neuron_parameter[206] <= 368'b11101010101010000010010000111100100100000001011001101010001101000111111101011001000000010000001000001001110010001001011111011110001110011111000111111010000000001011100000110000110110101100111001001000010000010000010001010011011101100110010110011010000000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011100000;
neuron_parameter[207] <= 368'b00011100001101010110100101100110011100010111001100100101000000111001101001101100001011011010000000000000010010010011010100000011111001010000101100011000001100011100100110101101001001100101000010100000000110101001101011001000100000010010101000100001111001000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110011110000;
neuron_parameter[208] <= 368'b10101001100010101100111110101010011111011010101010101000100010111010101010101110101110100010101010100010100010111010101010101010001010101010100011101010101010100010101010100010000110101010101010111110101010101011101010111010000110101010101000111110001000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100000000;
neuron_parameter[209] <= 368'b11111000001101011110101111100110011000011010000100101101011010010000000000101001101100001001101001111110000001010000100111011001010001100000100100101000000100100000100101100010010010011110100100101010100111000110100110001000100000000010101011010110111011010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100010000;
neuron_parameter[210] <= 368'b10100111110011101100010000011001000001101100111100011000010000100111111101101011100011110010011100000111111011001011000101000011111110101001111001000111001110100111010000000010011010011111001001101110000010100001001110011000010000111110000010001000100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100100000;
neuron_parameter[211] <= 368'b01110000101000100000001111100111111000011101010001100111101011010000000010111100000010001110101011001010011101010010100001001000101000001111101010011010111110001010101110101000010010101111100011101111110010100001111011011110001110101101011010001000111001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110100110000;
neuron_parameter[212] <= 368'b10100000100010110010101000011000000010101110100011001000110000100100010001110011010010001010001111101101111000001101111010001100100010000000000000000010000001010000001000001101001010100000010100100100001000001000001101100110101000101101011010010010100000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110101000000;
neuron_parameter[213] <= 368'b10011000101011101100111010101010111010110010101011101000101000111010101110101110100110101010101010101010110010011110101010101010101110001110101010101000101011001010101110101010001001101110101010101000101011101110101010111000101010101111001011101010100010110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110101010000;
neuron_parameter[214] <= 368'b00010110100001010010111100100010001110000010000001000101101100101011111100010110000001101101010000000001000110000011010010100000011110011100111111001101000010000111010110101011001100010111110010011010111110110001010110010101010111100001000110001010100101110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110101100000;
neuron_parameter[215] <= 368'b10000000110101000001001100000010001001100011000001000000010010011011010100101100100110100101111001100000100000010010000101000101010111011111000100111010110101110110111001011001110111101000110110000010110110000010010100100001010000100010101000110011010110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110101110000;
neuron_parameter[216] <= 368'b01101010000010010000000000011000100000000101000100001010101101001110111111011000100000100100101010101010100010101001011010100010000101111111000010001010110111001011101001110000100110001000111010011000000010010001110010111010111111000000110000001100001000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110000000;
neuron_parameter[217] <= 368'b00001101001010101110010010110110011110011100100110100011000001100000000010001011001100001000000011111011000101000101101010011000101001000000001010000000001000000100101000001100001101000000001100100000111000001010001110000000011000100001100000111011101110100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110010000;
neuron_parameter[218] <= 368'b10101011101010111000000010001001011011010010010000101000000100101101011011101011110000101110001010110110010110101101101101110111101110101110100100101010011000010000101110101110111000001011100000010010100000001111101001001100000000001110111100000000001011010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110100000;
neuron_parameter[219] <= 368'b11010010000101000000100011100100011100011001100010000101101011111001101101101110011101010100110111110010101110011110011011110100010000110001110101000100011010110010100000100010011000011111000000000001001111101110100111001001000000010111101001101101111011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110110110000;
neuron_parameter[220] <= 368'b11100101111011001000000010001000001011100010010100101000010101100111111101111000100010110010011000001000111010001011001101000010000011101001000000110001101001100011100001010010100000001011011011011111000000101010011010101010101000010001100000101101110011100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111000000;
neuron_parameter[221] <= 368'b00010010001100110111110100111011010110001100001000000011111010000010000000011001101010001010001001001110011000001011100001001100000001001011100010010000110001010111100110101110000111101000110110010101011000110000110000000000011101100101100010101000101011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111010000;
neuron_parameter[222] <= 368'b00100000110001010001110000001010100010101110101011101010110010110100010101110011010000101000000111101101101100001101100010001001101001000000101011000010001000001000001011001001001101000000000000100101001101100100000100001010101000101101011011110010100101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111100000;
neuron_parameter[223] <= 368'b10101110111110111010111010101010111010101010101010101010101110111011001000101010101110101010000010101010101010011010101010101010101010111010011110100010101011001011001010101010100010111010011111101010101011100000100110111010001000101001001011111000100110010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000110111110000;
neuron_parameter[224] <= 368'b00010000100000000100111011100011101100011010000000000100000010011001110010100110000101100100010101000000001110010010010101000000011110011100110101001111100110000010110110101001001000011101110010010110111110111001010110110100010111010001000000001010100001010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111000000000;
neuron_parameter[225] <= 368'b10100100100100001010000010110000100010110001001010110000110010101001000000000000101110001001100000101000110000010100010111001011110011111001000100101011111100101110111110001001100000101010000101001010110110010011010010111001001000001010111010000010001010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111000010000;
neuron_parameter[226] <= 368'b10101010111111100000010011000010100101000100001000011010001010110111100111011001010000110110000010010111011101001010011101011110000101011111000001001001010000000011100000110000110110010101101010001010111010010011010010110011011111000011110110111000000100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111000100000;
neuron_parameter[227] <= 368'b00000000101101001100100101100110111100010101001100100101001010110010001110111101001010011000100000000001000010000001010110000111110001010000001000100000001000011100010110001111011011100100000110100000101110111110011111001000000000111110101110100001101110000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111000110000;
neuron_parameter[228] <= 368'b10101001100010101010110010001011001010100010110010111000001110101101000010101010110000101110001110011110000010101100101101111101001110101110100101011000011000100100101001100100011100001111110000000100100101001111100001001000001000011110101011010000001011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001000000;
neuron_parameter[229] <= 368'b10010000001101000000111010100111111111010000100000100101100011011001101011001110001100101010111111111010101000011110011111110001101000101000110011001001001111100100101000101010011010101111000000010000111101110110100110101000001000110011101010111000111010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001010000;
neuron_parameter[230] <= 368'b00100111110011111000010000011000000010100110011101011010010100100111101101101011100011010010011000001111111011001011001001000010101010101001011001100001100011110111100000000010101010001011001001011110000011100110111110001100010000110010001010001000111000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001100000;
neuron_parameter[231] <= 368'b00010001001100010010001100000011000100010010000011010011111011100000000010010101011010001000001010001001001100000101100011001000100000010101010000010100110111010111110110101000000011101001010010010010111010110001111010010100110111110001100011001100110001100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111001110000;
neuron_parameter[232] <= 368'b00100011100010010111000000011001000000001000110011001000100001000100110011100010100011011011001000101101101000001001111010001110000000000001011011000101001001110000001000000000001111000000000100100100000000101000000101000010101000101111011110110001000100000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010000000;
neuron_parameter[233] <= 368'b11101101110110011000000000011001000001100110001100001000010000100111001001000011100000001101000000110111001000110101101100011101010100110110000100011010010000010111001110101011101011101010000100000101010001110100110001001000000000000101101001100000100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010010000;
neuron_parameter[234] <= 368'b00010110000001000010101001100110010110010010011001110111111111101000111001000110001101110100110101111011001011001000011011111010001010011010110100000101101010000001010111100001100100010111110010011011111011101111010000111100010111010001000101001100000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010100000;
neuron_parameter[235] <= 368'b11100101110010011000001000100100011000110101100010100000110010001010000100100000001110001000111101100000100000010011100101001101010111101111100110101011110101100100101001100001100110101100110100011001100110011010000010100001000001000110001000100001010100110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111010110000;
neuron_parameter[236] <= 368'b00100110100011100011000111000111001000110001001001011000101110100010100011111011010000110000101110100110100010101010000010110010000101001111110110001000101000001010101000010000100100101100101001011010011010010000110000100110010111000010010100001110000100010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011000000;
neuron_parameter[237] <= 368'b11010001011101001100101000010001110001010000101010100001000000011011101000111000001110000010100000000001100111100010000101000010001010111011110001100001101010011111110111100000111011011111010010001010100010111000000010001001001010101011101110001010001110110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011010000;
neuron_parameter[238] <= 368'b11101111110011111000110010011000000111100001011110101000000101101101000001001011111000101110000010110010011010111101111011111001000000111110100101101111011010110000011110101011101000101111100011001111101000000010001000011100000010001101001110100000111101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011100000;
neuron_parameter[239] <= 368'b01010010001100000000100101001000011100011000111000000101001001011001001100111100011111100000110001000001000001000010000101010000001010111010110101000101100010001011010101100010011010010111010000000000100000100000101001000000100010111011011100001000100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111011110000;
neuron_parameter[240] <= 368'b10101111101010101010010000011000000000100100010111111000100101100111101101101010100010010010011100001101111010001011001101000010110100011001100001001100001110100111100010000010110000111111001001001000000000100001000111000010011010110111000110101011100010000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100000000;
neuron_parameter[241] <= 368'b00010010000010110111111100001011110100000010000001010011101100000100000001010001111010001001101000001000011100010111100001001101110010010001101110110010111101001110101110001001001000101100010111111001011000110101011000010110111011000000000000001100010101100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100010000;
neuron_parameter[242] <= 368'b10100110100110001010000000101000111110100000101111101010011110101010111100010111100001111101001000100001100010000001100010101101100001000100000001101000100000011000000010001001001011101000110010101110001000100000001100000111010000101010001110000001011000010000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100100000;
neuron_parameter[243] <= 368'b10101001110101001001001000000100001011110011000000001000010100011011001000000100000101010100110001110000000000110100111100111001100000010000011110010100001010011100010110001101001100110111000000100110001100100000001100000010100000101000000111110011100011000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111100110000;
neuron_parameter[244] <= 368'b00010000000000100110111101100010011110000010101001000111001010011000111010000110110101101100100101100000000111010000010011100000001010011010111111100111100011100001000001100000001110011111111000010010110000111001010000010100010111011100000100000000000001110000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101000000;
neuron_parameter[245] <= 368'b00000000010000001000100100011000111001010001000010110100010000110010000100000000101010100000101111101000111001110100110011101011111010111011000000111101110100111110011100100010101001100010000110011101111100110000001010011000000010100001101011010000110010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101010000;
neuron_parameter[246] <= 368'b01101010010110101000010000011000100100000110001000101000101001001101111101001000100000110111001010101010110110101000101010000110000101001111000010001010100011001011101001100001100110101000111001001000100011011011100010111011111111000000110000000110001000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101100000;
neuron_parameter[247] <= 368'b00011010001001000000101101000110101010001011000000000101001010011000111000101100001011110010100000000001100111110010000101000011000010000001001000101100000010110101100010101100001011001001100110010110001001100111001101011010010010100010000111010100011101000000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111101110000;
neuron_parameter[248] <= 368'b00101110111000110000110101011001100010000100001100001010101010000110100011010001011001010111000110110011011100101101111010101010001000000110101110100101001010100100000101010011011000010101000001000000000010110000011010001000000100011000011000011001101000100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111110000000;
neuron_parameter[249] <= 368'b00100000111000000001101011101010111110111000001010101010101000001011101010101011001110101010101010001010101010000001100010101010101000001010101010101010101010101010101010101110101010001110101000100111001000100110101010100110001001000000001011111010110010100000000000000000000000000011111111110000000011111111110000000000000000000000000000000000001000000000111110010000;
neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;

            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
    else begin
        always @(negedge clk, negedge reset_n) begin
            if(~reset_n) begin
                neuron_parameter[0] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[1] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[2] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[3] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[4] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[5] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[6] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[7] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[8] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[9] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[10] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[11] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[12] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[13] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[14] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[15] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[16] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[17] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[18] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[19] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[20] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[21] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[22] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[23] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[24] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[25] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[26] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[27] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[28] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[29] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[30] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[31] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[32] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[33] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[34] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[35] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[36] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[37] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[38] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[39] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[40] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[41] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[42] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[43] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[44] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[45] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[46] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[47] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[48] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[49] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[50] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[51] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[52] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[53] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[54] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[55] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[56] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[57] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[58] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[59] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[60] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[61] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[62] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[63] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[64] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[65] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[66] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[67] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[68] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[69] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[70] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[71] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[72] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[73] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[74] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[75] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[76] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[77] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[78] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[79] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[80] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[81] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[82] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[83] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[84] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[85] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[86] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[87] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[88] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[89] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[90] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[91] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[92] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[93] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[94] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[95] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[96] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[97] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[98] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[99] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[100] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[101] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[102] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[103] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[104] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[105] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[106] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[107] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[108] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[109] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[110] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[111] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[112] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[113] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[114] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[115] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[116] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[117] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[118] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[119] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[120] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[121] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[122] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[123] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[124] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[125] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[126] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[127] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[128] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[129] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[130] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[131] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[132] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[133] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[134] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[135] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[136] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[137] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[138] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[139] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[140] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[141] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[142] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[143] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[144] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[145] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[146] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[147] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[148] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[149] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[150] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[151] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[152] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[153] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[154] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[155] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[156] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[157] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[158] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[159] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[160] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[161] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[162] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[163] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[164] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[165] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[166] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[167] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[168] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[169] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[170] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[171] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[172] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[173] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[174] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[175] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[176] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[177] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[178] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[179] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[180] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[181] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[182] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[183] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[184] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[185] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[186] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[187] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[188] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[189] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[190] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[191] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[192] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[193] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[194] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[195] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[196] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[197] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[198] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[199] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[200] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[201] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[202] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[203] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[204] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[205] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[206] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[207] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[208] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[209] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[210] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[211] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[212] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[213] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[214] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[215] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[216] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[217] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[218] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[219] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[220] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[221] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[222] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[223] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[224] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[225] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[226] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[227] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[228] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[229] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[230] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[231] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[232] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[233] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[234] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[235] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[236] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[237] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[238] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[239] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[240] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[241] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[242] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[243] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[244] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[245] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[246] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[247] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[248] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[249] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[250] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[251] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[252] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[253] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[254] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
                neuron_parameter[255] <= 368'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
            end
            else if(update_potential) begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i][111:103] <= potential_out[i];
            end
            else begin
                for(i = 0; i<256; i = i + 1) neuron_parameter[i] <= neuron_parameter[i];
            end
        end
    end
endgenerate

assign neuron_instructions[0] = 2'b00;
assign neuron_instructions[1] = 2'b01;
assign neuron_instructions[2] = 2'b00;
assign neuron_instructions[3] = 2'b01;
assign neuron_instructions[4] = 2'b00;
assign neuron_instructions[5] = 2'b01;
assign neuron_instructions[6] = 2'b00;
assign neuron_instructions[7] = 2'b01;
assign neuron_instructions[8] = 2'b00;
assign neuron_instructions[9] = 2'b01;
assign neuron_instructions[10] = 2'b00;
assign neuron_instructions[11] = 2'b01;
assign neuron_instructions[12] = 2'b00;
assign neuron_instructions[13] = 2'b01;
assign neuron_instructions[14] = 2'b00;
assign neuron_instructions[15] = 2'b01;
assign neuron_instructions[16] = 2'b00;
assign neuron_instructions[17] = 2'b01;
assign neuron_instructions[18] = 2'b00;
assign neuron_instructions[19] = 2'b01;
assign neuron_instructions[20] = 2'b00;
assign neuron_instructions[21] = 2'b01;
assign neuron_instructions[22] = 2'b00;
assign neuron_instructions[23] = 2'b01;
assign neuron_instructions[24] = 2'b00;
assign neuron_instructions[25] = 2'b01;
assign neuron_instructions[26] = 2'b00;
assign neuron_instructions[27] = 2'b01;
assign neuron_instructions[28] = 2'b00;
assign neuron_instructions[29] = 2'b01;
assign neuron_instructions[30] = 2'b00;
assign neuron_instructions[31] = 2'b01;
assign neuron_instructions[32] = 2'b00;
assign neuron_instructions[33] = 2'b01;
assign neuron_instructions[34] = 2'b00;
assign neuron_instructions[35] = 2'b01;
assign neuron_instructions[36] = 2'b00;
assign neuron_instructions[37] = 2'b01;
assign neuron_instructions[38] = 2'b00;
assign neuron_instructions[39] = 2'b01;
assign neuron_instructions[40] = 2'b00;
assign neuron_instructions[41] = 2'b01;
assign neuron_instructions[42] = 2'b00;
assign neuron_instructions[43] = 2'b01;
assign neuron_instructions[44] = 2'b00;
assign neuron_instructions[45] = 2'b01;
assign neuron_instructions[46] = 2'b00;
assign neuron_instructions[47] = 2'b01;
assign neuron_instructions[48] = 2'b00;
assign neuron_instructions[49] = 2'b01;
assign neuron_instructions[50] = 2'b00;
assign neuron_instructions[51] = 2'b01;
assign neuron_instructions[52] = 2'b00;
assign neuron_instructions[53] = 2'b01;
assign neuron_instructions[54] = 2'b00;
assign neuron_instructions[55] = 2'b01;
assign neuron_instructions[56] = 2'b00;
assign neuron_instructions[57] = 2'b01;
assign neuron_instructions[58] = 2'b00;
assign neuron_instructions[59] = 2'b01;
assign neuron_instructions[60] = 2'b00;
assign neuron_instructions[61] = 2'b01;
assign neuron_instructions[62] = 2'b00;
assign neuron_instructions[63] = 2'b01;
assign neuron_instructions[64] = 2'b00;
assign neuron_instructions[65] = 2'b01;
assign neuron_instructions[66] = 2'b00;
assign neuron_instructions[67] = 2'b01;
assign neuron_instructions[68] = 2'b00;
assign neuron_instructions[69] = 2'b01;
assign neuron_instructions[70] = 2'b00;
assign neuron_instructions[71] = 2'b01;
assign neuron_instructions[72] = 2'b00;
assign neuron_instructions[73] = 2'b01;
assign neuron_instructions[74] = 2'b00;
assign neuron_instructions[75] = 2'b01;
assign neuron_instructions[76] = 2'b00;
assign neuron_instructions[77] = 2'b01;
assign neuron_instructions[78] = 2'b00;
assign neuron_instructions[79] = 2'b01;
assign neuron_instructions[80] = 2'b00;
assign neuron_instructions[81] = 2'b01;
assign neuron_instructions[82] = 2'b00;
assign neuron_instructions[83] = 2'b01;
assign neuron_instructions[84] = 2'b00;
assign neuron_instructions[85] = 2'b01;
assign neuron_instructions[86] = 2'b00;
assign neuron_instructions[87] = 2'b01;
assign neuron_instructions[88] = 2'b00;
assign neuron_instructions[89] = 2'b01;
assign neuron_instructions[90] = 2'b00;
assign neuron_instructions[91] = 2'b01;
assign neuron_instructions[92] = 2'b00;
assign neuron_instructions[93] = 2'b01;
assign neuron_instructions[94] = 2'b00;
assign neuron_instructions[95] = 2'b01;
assign neuron_instructions[96] = 2'b00;
assign neuron_instructions[97] = 2'b01;
assign neuron_instructions[98] = 2'b00;
assign neuron_instructions[99] = 2'b01;
assign neuron_instructions[100] = 2'b00;
assign neuron_instructions[101] = 2'b01;
assign neuron_instructions[102] = 2'b00;
assign neuron_instructions[103] = 2'b01;
assign neuron_instructions[104] = 2'b00;
assign neuron_instructions[105] = 2'b01;
assign neuron_instructions[106] = 2'b00;
assign neuron_instructions[107] = 2'b01;
assign neuron_instructions[108] = 2'b00;
assign neuron_instructions[109] = 2'b01;
assign neuron_instructions[110] = 2'b00;
assign neuron_instructions[111] = 2'b01;
assign neuron_instructions[112] = 2'b00;
assign neuron_instructions[113] = 2'b01;
assign neuron_instructions[114] = 2'b00;
assign neuron_instructions[115] = 2'b01;
assign neuron_instructions[116] = 2'b00;
assign neuron_instructions[117] = 2'b01;
assign neuron_instructions[118] = 2'b00;
assign neuron_instructions[119] = 2'b01;
assign neuron_instructions[120] = 2'b00;
assign neuron_instructions[121] = 2'b01;
assign neuron_instructions[122] = 2'b00;
assign neuron_instructions[123] = 2'b01;
assign neuron_instructions[124] = 2'b00;
assign neuron_instructions[125] = 2'b01;
assign neuron_instructions[126] = 2'b00;
assign neuron_instructions[127] = 2'b01;
assign neuron_instructions[128] = 2'b00;
assign neuron_instructions[129] = 2'b01;
assign neuron_instructions[130] = 2'b00;
assign neuron_instructions[131] = 2'b01;
assign neuron_instructions[132] = 2'b00;
assign neuron_instructions[133] = 2'b01;
assign neuron_instructions[134] = 2'b00;
assign neuron_instructions[135] = 2'b01;
assign neuron_instructions[136] = 2'b00;
assign neuron_instructions[137] = 2'b01;
assign neuron_instructions[138] = 2'b00;
assign neuron_instructions[139] = 2'b01;
assign neuron_instructions[140] = 2'b00;
assign neuron_instructions[141] = 2'b01;
assign neuron_instructions[142] = 2'b00;
assign neuron_instructions[143] = 2'b01;
assign neuron_instructions[144] = 2'b00;
assign neuron_instructions[145] = 2'b01;
assign neuron_instructions[146] = 2'b00;
assign neuron_instructions[147] = 2'b01;
assign neuron_instructions[148] = 2'b00;
assign neuron_instructions[149] = 2'b01;
assign neuron_instructions[150] = 2'b00;
assign neuron_instructions[151] = 2'b01;
assign neuron_instructions[152] = 2'b00;
assign neuron_instructions[153] = 2'b01;
assign neuron_instructions[154] = 2'b00;
assign neuron_instructions[155] = 2'b01;
assign neuron_instructions[156] = 2'b00;
assign neuron_instructions[157] = 2'b01;
assign neuron_instructions[158] = 2'b00;
assign neuron_instructions[159] = 2'b01;
assign neuron_instructions[160] = 2'b00;
assign neuron_instructions[161] = 2'b01;
assign neuron_instructions[162] = 2'b00;
assign neuron_instructions[163] = 2'b01;
assign neuron_instructions[164] = 2'b00;
assign neuron_instructions[165] = 2'b01;
assign neuron_instructions[166] = 2'b00;
assign neuron_instructions[167] = 2'b01;
assign neuron_instructions[168] = 2'b00;
assign neuron_instructions[169] = 2'b01;
assign neuron_instructions[170] = 2'b00;
assign neuron_instructions[171] = 2'b01;
assign neuron_instructions[172] = 2'b00;
assign neuron_instructions[173] = 2'b01;
assign neuron_instructions[174] = 2'b00;
assign neuron_instructions[175] = 2'b01;
assign neuron_instructions[176] = 2'b00;
assign neuron_instructions[177] = 2'b01;
assign neuron_instructions[178] = 2'b00;
assign neuron_instructions[179] = 2'b01;
assign neuron_instructions[180] = 2'b00;
assign neuron_instructions[181] = 2'b01;
assign neuron_instructions[182] = 2'b00;
assign neuron_instructions[183] = 2'b01;
assign neuron_instructions[184] = 2'b00;
assign neuron_instructions[185] = 2'b01;
assign neuron_instructions[186] = 2'b00;
assign neuron_instructions[187] = 2'b01;
assign neuron_instructions[188] = 2'b00;
assign neuron_instructions[189] = 2'b01;
assign neuron_instructions[190] = 2'b00;
assign neuron_instructions[191] = 2'b01;
assign neuron_instructions[192] = 2'b00;
assign neuron_instructions[193] = 2'b01;
assign neuron_instructions[194] = 2'b00;
assign neuron_instructions[195] = 2'b01;
assign neuron_instructions[196] = 2'b00;
assign neuron_instructions[197] = 2'b01;
assign neuron_instructions[198] = 2'b00;
assign neuron_instructions[199] = 2'b01;
assign neuron_instructions[200] = 2'b00;
assign neuron_instructions[201] = 2'b01;
assign neuron_instructions[202] = 2'b00;
assign neuron_instructions[203] = 2'b01;
assign neuron_instructions[204] = 2'b00;
assign neuron_instructions[205] = 2'b01;
assign neuron_instructions[206] = 2'b00;
assign neuron_instructions[207] = 2'b01;
assign neuron_instructions[208] = 2'b00;
assign neuron_instructions[209] = 2'b01;
assign neuron_instructions[210] = 2'b00;
assign neuron_instructions[211] = 2'b01;
assign neuron_instructions[212] = 2'b00;
assign neuron_instructions[213] = 2'b01;
assign neuron_instructions[214] = 2'b00;
assign neuron_instructions[215] = 2'b01;
assign neuron_instructions[216] = 2'b00;
assign neuron_instructions[217] = 2'b01;
assign neuron_instructions[218] = 2'b00;
assign neuron_instructions[219] = 2'b01;
assign neuron_instructions[220] = 2'b00;
assign neuron_instructions[221] = 2'b01;
assign neuron_instructions[222] = 2'b00;
assign neuron_instructions[223] = 2'b01;
assign neuron_instructions[224] = 2'b00;
assign neuron_instructions[225] = 2'b01;
assign neuron_instructions[226] = 2'b00;
assign neuron_instructions[227] = 2'b01;
assign neuron_instructions[228] = 2'b00;
assign neuron_instructions[229] = 2'b01;
assign neuron_instructions[230] = 2'b00;
assign neuron_instructions[231] = 2'b01;
assign neuron_instructions[232] = 2'b00;
assign neuron_instructions[233] = 2'b01;
assign neuron_instructions[234] = 2'b00;
assign neuron_instructions[235] = 2'b01;
assign neuron_instructions[236] = 2'b00;
assign neuron_instructions[237] = 2'b01;
assign neuron_instructions[238] = 2'b00;
assign neuron_instructions[239] = 2'b01;
assign neuron_instructions[240] = 2'b00;
assign neuron_instructions[241] = 2'b01;
assign neuron_instructions[242] = 2'b00;
assign neuron_instructions[243] = 2'b01;
assign neuron_instructions[244] = 2'b00;
assign neuron_instructions[245] = 2'b01;
assign neuron_instructions[246] = 2'b00;
assign neuron_instructions[247] = 2'b01;
assign neuron_instructions[248] = 2'b00;
assign neuron_instructions[249] = 2'b01;
assign neuron_instructions[250] = 2'b00;
assign neuron_instructions[251] = 2'b01;
assign neuron_instructions[252] = 2'b00;
assign neuron_instructions[253] = 2'b01;
assign neuron_instructions[254] = 2'b00;
assign neuron_instructions[255] = 2'b01;
endmodule

